magic
tech sky130B
timestamp 1647929098
<< nwell >>
rect 3011 -200 3139 -170
rect 2975 -327 3139 -200
<< metal1 >>
rect 5336 5207 5409 5223
rect 5336 3109 5344 5207
rect 5397 3109 5409 5207
rect 2925 3093 2975 3108
rect 2925 3052 2932 3093
rect 2969 3052 2975 3093
rect 2925 3040 2975 3052
rect 4728 3092 4774 3098
rect 5336 3093 5409 3109
rect 4728 3053 4734 3092
rect 4769 3053 4774 3092
rect 2935 3009 2965 3040
rect 4728 3029 4774 3053
rect 5356 3030 5381 3093
rect 5166 -187 5191 -170
rect 3009 -228 5191 -187
rect -326 -1913 -214 -1907
rect -326 -1947 -319 -1913
rect -277 -1947 -214 -1913
rect -326 -1953 -214 -1947
rect 3009 -2070 3051 -228
rect 2972 -2095 3051 -2070
<< via1 >>
rect 5344 3109 5397 5207
rect 2932 3052 2969 3093
rect 4734 3053 4769 3092
rect -319 -1947 -277 -1913
<< metal2 >>
rect 5336 5207 5409 5223
rect 5336 3109 5344 5207
rect 5397 3109 5409 5207
rect 2925 3093 2975 3108
rect 2925 3052 2932 3093
rect 2969 3052 2975 3093
rect 2925 3040 2975 3052
rect 4728 3092 4775 3098
rect 5336 3093 5409 3109
rect 4728 3053 4734 3092
rect 4769 3053 4775 3092
rect 4728 3048 4775 3053
rect -328 -162 -266 -156
rect -328 -198 -323 -162
rect -272 -175 -266 -162
rect -272 -190 -215 -175
rect -272 -198 -266 -190
rect -328 -207 -266 -198
rect -326 -1913 -269 -1907
rect -326 -1948 -320 -1913
rect -277 -1948 -269 -1913
rect -326 -1954 -269 -1948
<< via2 >>
rect 5344 3109 5397 5207
rect 2932 3052 2969 3093
rect 4734 3053 4769 3085
rect -323 -198 -272 -162
rect -320 -1947 -319 -1913
rect -319 -1947 -277 -1913
rect -320 -1948 -277 -1947
<< metal3 >>
rect 5650 5236 30750 15050
rect 5319 5207 30750 5236
rect 2925 3093 2975 3108
rect 2925 3052 2932 3093
rect 2969 3052 2975 3093
rect 2925 3040 2975 3052
rect 4716 3085 4785 3127
rect 5319 3109 5344 5207
rect 5397 3109 30750 5207
rect 5319 3093 30750 3109
rect 4716 3053 4734 3085
rect 4769 3053 4785 3085
rect 4716 3042 4785 3053
rect -331 -162 -266 -153
rect -331 -198 -323 -162
rect -272 -198 -266 -162
rect -331 -212 -266 -198
rect -327 -1913 -269 -1907
rect -327 -1948 -320 -1913
rect -277 -1948 -269 -1913
rect -327 -1954 -269 -1948
rect 5650 -10050 30750 3093
<< via3 >>
rect 2932 3052 2969 3093
rect 4734 3053 4769 3085
rect -323 -198 -272 -162
rect -320 -1948 -277 -1913
<< mimcap >>
rect 5700 14000 30700 15000
rect 5700 12000 6000 14000
rect 30000 12000 30700 14000
rect 5700 -7000 30700 12000
rect 5700 -9000 6000 -7000
rect 30000 -9000 30700 -7000
rect 5700 -10000 30700 -9000
<< mimcapcontact >>
rect 6000 12000 30000 14000
rect 6000 -9000 30000 -7000
<< metal4 >>
rect 5660 14000 30760 15050
rect 5660 12000 6000 14000
rect 30000 12000 30760 14000
rect 5660 5237 30760 12000
rect 2925 3098 2975 3108
rect 4427 3098 30760 5237
rect 2565 3093 30760 3098
rect 2565 3052 2932 3093
rect 2969 3085 30760 3093
rect 2969 3053 4734 3085
rect 4769 3053 30760 3085
rect 2969 3052 30760 3053
rect 2565 3048 30760 3052
rect 2925 3040 2975 3048
rect -331 -162 -266 -153
rect -331 -198 -323 -162
rect -272 -198 -266 -162
rect -331 -212 -266 -198
rect -326 -1913 -269 -212
rect -326 -1948 -320 -1913
rect -277 -1948 -269 -1913
rect -326 -1953 -269 -1948
rect 5660 -7000 30760 3048
rect 5660 -9000 6000 -7000
rect 30000 -9000 30760 -7000
rect 5660 -10050 30760 -9000
use 1T1R_16x16  1T1R_16x16_0 ~/Desktop/cmos_reram
timestamp 1647888104
transform 1 0 -225 0 1 -195
box 0 -35 3200 3205
use col_driver_1x2  col_driver_1x2_0 ~/Desktop/cmos_reram
timestamp 1647923593
transform 1 0 -225 0 1 -2485
box 0 0 400 2305
use col_driver_1x2  col_driver_1x2_1
timestamp 1647923593
transform 1 0 175 0 1 -2485
box 0 0 400 2305
use col_driver_1x2  col_driver_1x2_2
timestamp 1647923593
transform 1 0 575 0 1 -2485
box 0 0 400 2305
use col_driver_1x2  col_driver_1x2_3
timestamp 1647923593
transform 1 0 975 0 1 -2485
box 0 0 400 2305
use col_driver_1x2  col_driver_1x2_4
timestamp 1647923593
transform 1 0 1375 0 1 -2485
box 0 0 400 2305
use col_driver_1x2  col_driver_1x2_5
timestamp 1647923593
transform 1 0 1775 0 1 -2485
box 0 0 400 2305
use col_driver_1x2  col_driver_1x2_6
timestamp 1647923593
transform 1 0 2175 0 1 -2485
box 0 0 400 2305
use col_driver_1x2  col_driver_1x2_7
timestamp 1647923593
transform 1 0 2575 0 1 -2485
box 0 0 400 2305
use row_driver_2x1  row_driver_2x1_0 ~/Desktop/cmos_reram
timestamp 1647923593
transform 1 0 3041 0 1 2605
box -66 24 2445 425
use row_driver_2x1  row_driver_2x1_1
timestamp 1647923593
transform 1 0 3041 0 1 -195
box -66 24 2445 425
use row_driver_2x1  row_driver_2x1_2
timestamp 1647923593
transform 1 0 3041 0 1 205
box -66 24 2445 425
use row_driver_2x1  row_driver_2x1_3
timestamp 1647923593
transform 1 0 3041 0 1 605
box -66 24 2445 425
use row_driver_2x1  row_driver_2x1_4
timestamp 1647923593
transform 1 0 3041 0 1 1005
box -66 24 2445 425
use row_driver_2x1  row_driver_2x1_5
timestamp 1647923593
transform 1 0 3041 0 1 1405
box -66 24 2445 425
use row_driver_2x1  row_driver_2x1_6
timestamp 1647923593
transform 1 0 3041 0 1 1805
box -66 24 2445 425
use row_driver_2x1  row_driver_2x1_7
timestamp 1647923593
transform 1 0 3041 0 1 2205
box -66 24 2445 425
<< end >>
