VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO col_driver
  CLASS BLOCK ;
  FOREIGN col_driver ;
  ORIGIN 0.300 19.340 ;
  SIZE 2.000 BY 23.050 ;
  PIN Vgnc
    ANTENNAGATEAREA 1.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 -11.990 1.700 -11.590 ;
        RECT 1.300 -12.540 1.600 -11.990 ;
        RECT 1.200 -12.940 1.700 -12.540 ;
      LAYER mcon ;
        RECT 1.300 -11.940 1.600 -11.640 ;
        RECT 1.300 -12.890 1.600 -12.590 ;
      LAYER met1 ;
        RECT 1.200 -11.640 1.700 -11.590 ;
        RECT -0.300 -11.940 1.700 -11.640 ;
        RECT 1.200 -11.990 1.700 -11.940 ;
        RECT 1.200 -12.590 1.700 -12.540 ;
        RECT -0.300 -12.890 1.700 -12.590 ;
        RECT 1.200 -12.940 1.700 -12.890 ;
    END
  END Vgnc
  PIN Vref
    ANTENNADIFFAREA 1.350000 ;
    PORT
      LAYER li1 ;
        RECT -0.130 -15.490 1.000 -15.140 ;
        RECT -0.130 -17.040 0.040 -15.490 ;
        RECT -0.130 -17.390 1.000 -17.040 ;
        RECT -0.130 -18.940 0.040 -17.390 ;
        RECT -0.130 -19.290 1.000 -18.940 ;
      LAYER mcon ;
        RECT 0.200 -15.440 0.900 -15.190 ;
        RECT 0.200 -17.340 0.900 -17.090 ;
        RECT 0.200 -19.240 0.900 -18.990 ;
      LAYER met1 ;
        RECT 0.060 -15.190 1.000 -15.130 ;
        RECT -0.300 -15.440 1.700 -15.190 ;
        RECT 0.060 -15.490 1.000 -15.440 ;
        RECT 0.060 -17.090 1.000 -17.030 ;
        RECT -0.300 -17.340 1.700 -17.090 ;
        RECT 0.060 -17.390 1.000 -17.340 ;
        RECT 0.060 -18.990 1.000 -18.930 ;
        RECT -0.300 -19.240 1.700 -18.990 ;
        RECT 0.060 -19.290 1.000 -19.240 ;
    END
  END Vref
  PIN Vgpc
    ANTENNAGATEAREA 2.500000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 -2.540 1.700 -2.140 ;
        RECT 1.300 -3.090 1.600 -2.540 ;
        RECT 1.200 -3.490 1.700 -3.090 ;
        RECT 1.300 -4.040 1.600 -3.490 ;
        RECT 1.200 -4.440 1.700 -4.040 ;
        RECT 1.300 -4.990 1.600 -4.440 ;
        RECT 1.200 -5.390 1.700 -4.990 ;
        RECT 1.300 -5.940 1.600 -5.390 ;
        RECT 1.200 -6.340 1.700 -5.940 ;
      LAYER mcon ;
        RECT 1.300 -2.490 1.600 -2.190 ;
        RECT 1.300 -3.440 1.600 -3.140 ;
        RECT 1.300 -4.390 1.600 -4.090 ;
        RECT 1.300 -5.340 1.600 -5.040 ;
        RECT 1.300 -6.290 1.600 -5.990 ;
      LAYER met1 ;
        RECT 1.200 -2.190 1.700 -2.140 ;
        RECT -0.300 -2.490 1.700 -2.190 ;
        RECT 1.200 -2.540 1.700 -2.490 ;
        RECT 1.200 -3.490 1.700 -3.090 ;
        RECT 1.200 -4.440 1.700 -4.040 ;
        RECT 1.200 -5.390 1.700 -4.990 ;
        RECT 1.200 -6.340 1.700 -5.940 ;
    END
  END Vgpc
  PIN SWc_minus
    ANTENNAGATEAREA 2.500000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 -15.040 1.700 -14.640 ;
        RECT 1.200 -15.990 1.700 -15.590 ;
        RECT 1.200 -16.940 1.700 -16.540 ;
        RECT 1.200 -17.890 1.700 -17.490 ;
        RECT 1.200 -18.840 1.700 -18.440 ;
      LAYER mcon ;
        RECT 1.300 -14.990 1.600 -14.690 ;
        RECT 1.300 -15.940 1.600 -15.640 ;
        RECT 1.300 -16.890 1.600 -16.590 ;
        RECT 1.300 -17.840 1.600 -17.540 ;
        RECT 1.300 -18.790 1.600 -18.490 ;
      LAYER met1 ;
        RECT 1.200 -15.040 1.700 -14.640 ;
        RECT 1.200 -15.990 1.700 -15.590 ;
        RECT 1.200 -16.940 1.700 -16.540 ;
        RECT 1.200 -17.890 1.700 -17.490 ;
        RECT 1.200 -18.840 1.700 -18.440 ;
      LAYER via ;
        RECT 1.300 -14.990 1.600 -14.690 ;
        RECT 1.300 -15.940 1.600 -15.640 ;
        RECT 1.300 -16.890 1.600 -16.590 ;
        RECT 1.300 -17.840 1.600 -17.540 ;
        RECT 1.300 -18.790 1.600 -18.490 ;
      LAYER met2 ;
        RECT 1.200 -15.040 1.700 -14.640 ;
        RECT 1.350 -15.590 1.550 -15.040 ;
        RECT 1.200 -15.990 1.700 -15.590 ;
        RECT 1.350 -16.540 1.550 -15.990 ;
        RECT 1.200 -16.940 1.700 -16.540 ;
        RECT 1.350 -17.490 1.550 -16.940 ;
        RECT 1.200 -17.890 1.700 -17.490 ;
        RECT 1.350 -18.440 1.550 -17.890 ;
        RECT 1.200 -18.840 1.700 -18.440 ;
        RECT 1.350 -19.340 1.550 -18.840 ;
    END
  END SWc_minus
  PIN SWref
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 -9.140 1.700 -8.740 ;
        RECT 1.200 -10.090 1.700 -9.690 ;
        RECT 1.200 -11.040 1.700 -10.640 ;
      LAYER mcon ;
        RECT 1.300 -9.090 1.600 -8.790 ;
        RECT 1.300 -10.040 1.600 -9.740 ;
        RECT 1.300 -10.990 1.600 -10.690 ;
      LAYER met1 ;
        RECT 1.200 -9.140 1.700 -8.740 ;
        RECT 1.200 -10.090 1.700 -9.690 ;
        RECT 1.200 -11.040 1.700 -10.640 ;
      LAYER via ;
        RECT 1.300 -9.090 1.600 -8.790 ;
        RECT 1.300 -10.040 1.600 -9.740 ;
        RECT 1.300 -10.990 1.600 -10.690 ;
      LAYER met2 ;
        RECT 1.200 -9.140 1.700 -8.740 ;
        RECT 1.200 -10.090 1.700 -9.690 ;
        RECT 1.200 -11.040 1.700 -10.640 ;
      LAYER via2 ;
        RECT 1.300 -9.090 1.600 -8.790 ;
        RECT 1.300 -10.040 1.600 -9.740 ;
        RECT 1.300 -10.990 1.600 -10.690 ;
      LAYER met3 ;
        RECT 1.200 -9.190 1.700 -8.690 ;
        RECT 1.300 -9.640 1.600 -9.190 ;
        RECT 1.200 -10.140 1.700 -9.640 ;
        RECT 1.300 -10.590 1.600 -10.140 ;
        RECT 1.200 -11.090 1.700 -10.590 ;
        RECT 1.300 -19.340 1.600 -11.090 ;
    END
  END SWref
  PIN SWc_plus
    ANTENNAGATEAREA 2.500000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 2.210 1.700 2.610 ;
        RECT 1.200 1.260 1.700 1.660 ;
        RECT 1.200 0.310 1.700 0.710 ;
        RECT 1.200 -0.640 1.700 -0.240 ;
        RECT 1.200 -1.590 1.700 -1.190 ;
      LAYER mcon ;
        RECT 1.300 2.260 1.600 2.560 ;
        RECT 1.300 1.310 1.600 1.610 ;
        RECT 1.300 0.360 1.600 0.660 ;
        RECT 1.300 -0.590 1.600 -0.290 ;
        RECT 1.300 -1.540 1.600 -1.240 ;
      LAYER met1 ;
        RECT 1.200 2.210 1.700 2.610 ;
        RECT 1.200 1.260 1.700 1.660 ;
        RECT 1.200 0.310 1.700 0.710 ;
        RECT 1.200 -0.640 1.700 -0.240 ;
        RECT 1.200 -1.590 1.700 -1.190 ;
      LAYER via ;
        RECT 1.300 2.260 1.600 2.560 ;
        RECT 1.300 1.310 1.600 1.610 ;
        RECT 1.300 0.360 1.600 0.660 ;
        RECT 1.300 -0.590 1.600 -0.290 ;
        RECT 1.300 -1.540 1.600 -1.240 ;
      LAYER met2 ;
        RECT 1.200 2.210 1.700 2.610 ;
        RECT 1.200 1.260 1.700 1.660 ;
        RECT 1.200 0.310 1.700 0.710 ;
        RECT 1.200 -0.640 1.700 -0.240 ;
        RECT 1.200 -1.590 1.700 -1.190 ;
      LAYER via2 ;
        RECT 1.300 2.260 1.600 2.560 ;
        RECT 1.300 1.310 1.600 1.610 ;
        RECT 1.300 0.360 1.600 0.660 ;
        RECT 1.300 -0.590 1.600 -0.290 ;
        RECT 1.300 -1.540 1.600 -1.240 ;
      LAYER met3 ;
        RECT 1.200 2.160 1.700 2.660 ;
        RECT 1.200 1.210 1.700 1.710 ;
        RECT 1.200 0.260 1.700 0.760 ;
        RECT 1.200 -0.690 1.700 -0.190 ;
        RECT 1.200 -1.640 1.700 -1.140 ;
      LAYER via3 ;
        RECT 1.290 2.250 1.610 2.570 ;
        RECT 1.290 1.300 1.610 1.620 ;
        RECT 1.290 0.350 1.610 0.670 ;
        RECT 1.290 -0.600 1.610 -0.280 ;
        RECT 1.290 -1.550 1.610 -1.230 ;
      LAYER met4 ;
        RECT 1.200 2.210 1.700 2.610 ;
        RECT 1.300 1.660 1.600 2.210 ;
        RECT 1.200 1.260 1.700 1.660 ;
        RECT 1.300 0.710 1.600 1.260 ;
        RECT 1.200 0.310 1.700 0.710 ;
        RECT 1.300 -0.240 1.600 0.310 ;
        RECT 1.200 -0.640 1.700 -0.240 ;
        RECT 1.300 -1.190 1.600 -0.640 ;
        RECT 1.200 -1.590 1.700 -1.190 ;
        RECT 1.300 -2.140 1.600 -1.590 ;
        RECT 1.200 -2.540 1.700 -2.140 ;
        RECT 1.300 -3.090 1.600 -2.540 ;
        RECT 1.200 -3.490 1.700 -3.090 ;
        RECT 1.300 -4.040 1.600 -3.490 ;
        RECT 1.200 -4.440 1.700 -4.040 ;
        RECT 1.300 -4.990 1.600 -4.440 ;
        RECT 1.200 -5.390 1.700 -4.990 ;
        RECT 1.300 -5.940 1.600 -5.390 ;
        RECT 1.200 -6.340 1.700 -5.940 ;
        RECT 1.300 -19.340 1.600 -6.340 ;
    END
  END SWc_plus
  PIN Vc_minus
    ANTENNADIFFAREA 0.450000 ;
    PORT
      LAYER li1 ;
        RECT 0.210 -12.440 1.000 -12.090 ;
      LAYER mcon ;
        RECT 0.210 -12.390 0.900 -12.140 ;
      LAYER met1 ;
        RECT -0.150 -12.140 1.000 -12.090 ;
        RECT -0.300 -12.390 1.700 -12.140 ;
        RECT -0.150 -12.440 1.000 -12.390 ;
    END
  END Vc_minus
  PIN Vc_plus
    ANTENNADIFFAREA 1.350000 ;
    PORT
      LAYER li1 ;
        RECT 0.210 -2.990 1.000 -2.640 ;
        RECT 0.210 -4.890 1.000 -4.540 ;
        RECT 0.150 -6.790 1.000 -6.440 ;
      LAYER mcon ;
        RECT 0.250 -2.940 0.900 -2.690 ;
        RECT 0.250 -4.840 0.900 -4.590 ;
        RECT 0.250 -6.740 0.900 -6.490 ;
      LAYER met1 ;
        RECT 0.150 -2.690 1.000 -2.640 ;
        RECT -0.300 -2.940 1.700 -2.690 ;
        RECT -0.150 -4.590 0.000 -2.940 ;
        RECT 0.150 -2.990 1.000 -2.940 ;
        RECT 0.150 -4.590 1.000 -4.540 ;
        RECT -0.300 -4.840 1.700 -4.590 ;
        RECT -0.150 -6.490 0.000 -4.840 ;
        RECT 0.150 -4.890 1.000 -4.840 ;
        RECT 0.150 -6.490 1.000 -6.440 ;
        RECT -0.300 -6.740 1.700 -6.490 ;
        RECT 0.150 -6.790 1.000 -6.740 ;
    END
  END Vc_plus
  PIN vssd1
    ANTENNADIFFAREA 0.700000 ;
    PORT
      LAYER li1 ;
        RECT 0.210 -14.020 1.000 -13.560 ;
      LAYER mcon ;
        RECT 0.210 -13.980 0.900 -13.600 ;
      LAYER met1 ;
        RECT -0.300 -14.020 1.700 -13.560 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 0.700000 ;
    PORT
      LAYER nwell ;
        RECT -0.300 -7.890 1.700 3.510 ;
      LAYER li1 ;
        RECT 0.100 -7.490 1.000 -6.990 ;
      LAYER mcon ;
        RECT 0.200 -7.390 0.900 -7.090 ;
      LAYER met1 ;
        RECT -0.300 -7.440 1.700 -7.040 ;
    END
  END vccd1
  OBS
      LAYER li1 ;
        RECT 0.150 2.710 1.000 3.060 ;
        RECT -0.130 2.110 0.040 2.530 ;
        RECT -0.130 1.760 1.000 2.110 ;
        RECT -0.130 0.210 0.040 1.760 ;
        RECT 0.210 0.810 1.000 1.160 ;
        RECT -0.130 -0.140 1.000 0.210 ;
        RECT -0.130 -1.690 0.040 -0.140 ;
        RECT 0.210 -1.090 1.000 -0.740 ;
        RECT -0.130 -2.040 1.000 -1.690 ;
        RECT -0.130 -3.590 0.040 -2.040 ;
        RECT -0.130 -3.940 1.000 -3.590 ;
        RECT -0.130 -5.490 0.040 -3.940 ;
        RECT -0.130 -5.840 1.000 -5.490 ;
        RECT -0.130 -9.240 0.040 -8.240 ;
        RECT 0.210 -8.640 1.000 -8.290 ;
        RECT -0.130 -9.590 1.000 -9.240 ;
        RECT -0.130 -11.140 0.040 -9.590 ;
        RECT 0.210 -10.540 1.000 -10.190 ;
        RECT -0.130 -11.490 1.000 -11.140 ;
        RECT -0.130 -13.040 0.040 -11.490 ;
        RECT -0.130 -13.390 1.000 -13.040 ;
        RECT 0.100 -14.540 1.000 -14.190 ;
        RECT 0.210 -16.440 1.000 -16.090 ;
        RECT 0.210 -18.340 1.000 -17.990 ;
      LAYER mcon ;
        RECT 0.250 2.760 0.900 3.010 ;
        RECT 0.250 0.860 0.900 1.110 ;
        RECT 0.250 -1.040 0.900 -0.790 ;
        RECT 0.250 -8.590 0.900 -8.340 ;
        RECT 0.250 -10.490 0.900 -10.240 ;
        RECT 0.250 -14.490 0.900 -14.240 ;
        RECT 0.250 -16.390 0.900 -16.140 ;
        RECT 0.250 -18.290 0.900 -18.040 ;
      LAYER met1 ;
        RECT -0.250 3.510 0.660 3.710 ;
        RECT 0.460 3.060 0.660 3.510 ;
        RECT 0.150 2.710 1.000 3.060 ;
        RECT 0.150 0.810 1.000 1.160 ;
        RECT 0.150 -1.090 1.000 -0.740 ;
        RECT 0.150 -8.640 1.000 -8.290 ;
        RECT 0.150 -10.540 1.000 -10.190 ;
        RECT 0.150 -14.540 1.000 -14.190 ;
        RECT 0.150 -16.440 1.000 -16.090 ;
        RECT 0.150 -18.340 1.000 -17.990 ;
      LAYER via ;
        RECT 0.250 2.710 0.900 3.060 ;
        RECT 0.250 0.810 0.900 1.160 ;
        RECT 0.250 -1.090 0.900 -0.740 ;
        RECT 0.250 -8.640 0.900 -8.290 ;
        RECT 0.250 -10.540 0.900 -10.190 ;
        RECT 0.250 -14.540 0.900 -14.190 ;
        RECT 0.250 -16.440 0.900 -16.090 ;
        RECT 0.250 -18.340 0.900 -17.990 ;
      LAYER met2 ;
        RECT -0.150 2.710 1.000 3.060 ;
        RECT -0.150 1.160 0.050 2.710 ;
        RECT -0.150 0.810 1.000 1.160 ;
        RECT -0.150 -0.740 0.050 0.810 ;
        RECT -0.150 -1.090 1.000 -0.740 ;
        RECT -0.150 -8.290 0.050 -1.090 ;
        RECT -0.150 -8.640 1.000 -8.290 ;
        RECT -0.150 -10.190 0.050 -8.640 ;
        RECT -0.150 -10.540 1.000 -10.190 ;
        RECT -0.150 -14.190 0.050 -10.540 ;
        RECT -0.150 -14.540 1.000 -14.190 ;
        RECT -0.150 -16.090 0.050 -14.540 ;
        RECT -0.150 -16.440 1.000 -16.090 ;
        RECT -0.150 -17.990 0.050 -16.440 ;
        RECT -0.150 -18.340 1.000 -17.990 ;
        RECT -0.150 -19.290 0.050 -18.930 ;
  END
END col_driver
END LIBRARY

