magic
tech sky130B
timestamp 1647923593
use col_driver  col_driver_0
timestamp 1647920282
transform 1 0 30 0 1 1934
box -30 -1934 170 371
use col_driver  col_driver_1
timestamp 1647920282
transform 1 0 230 0 1 1934
box -30 -1934 170 371
<< end >>
