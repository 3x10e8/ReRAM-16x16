magic
tech sky130B
timestamp 1647720169
<< metal1 >>
rect -25 -15 15 25
<< reram >>
rect -20 -10 10 20
<< metal2 >>
rect -25 20 15 25
rect -25 -10 -20 20
rect 10 -10 15 20
rect -25 -15 15 -10
<< end >>
