magic
tech sky130A
magscale 1 2
timestamp 1609532432
<< pwell >>
rect -2521 -827 2521 827
<< mvnmos >>
rect -2293 -569 -2093 631
rect -2035 -569 -1835 631
rect -1777 -569 -1577 631
rect -1519 -569 -1319 631
rect -1261 -569 -1061 631
rect -1003 -569 -803 631
rect -745 -569 -545 631
rect -487 -569 -287 631
rect -229 -569 -29 631
rect 29 -569 229 631
rect 287 -569 487 631
rect 545 -569 745 631
rect 803 -569 1003 631
rect 1061 -569 1261 631
rect 1319 -569 1519 631
rect 1577 -569 1777 631
rect 1835 -569 2035 631
rect 2093 -569 2293 631
<< mvndiff >>
rect -2351 619 -2293 631
rect -2351 -557 -2339 619
rect -2305 -557 -2293 619
rect -2351 -569 -2293 -557
rect -2093 619 -2035 631
rect -2093 -557 -2081 619
rect -2047 -557 -2035 619
rect -2093 -569 -2035 -557
rect -1835 619 -1777 631
rect -1835 -557 -1823 619
rect -1789 -557 -1777 619
rect -1835 -569 -1777 -557
rect -1577 619 -1519 631
rect -1577 -557 -1565 619
rect -1531 -557 -1519 619
rect -1577 -569 -1519 -557
rect -1319 619 -1261 631
rect -1319 -557 -1307 619
rect -1273 -557 -1261 619
rect -1319 -569 -1261 -557
rect -1061 619 -1003 631
rect -1061 -557 -1049 619
rect -1015 -557 -1003 619
rect -1061 -569 -1003 -557
rect -803 619 -745 631
rect -803 -557 -791 619
rect -757 -557 -745 619
rect -803 -569 -745 -557
rect -545 619 -487 631
rect -545 -557 -533 619
rect -499 -557 -487 619
rect -545 -569 -487 -557
rect -287 619 -229 631
rect -287 -557 -275 619
rect -241 -557 -229 619
rect -287 -569 -229 -557
rect -29 619 29 631
rect -29 -557 -17 619
rect 17 -557 29 619
rect -29 -569 29 -557
rect 229 619 287 631
rect 229 -557 241 619
rect 275 -557 287 619
rect 229 -569 287 -557
rect 487 619 545 631
rect 487 -557 499 619
rect 533 -557 545 619
rect 487 -569 545 -557
rect 745 619 803 631
rect 745 -557 757 619
rect 791 -557 803 619
rect 745 -569 803 -557
rect 1003 619 1061 631
rect 1003 -557 1015 619
rect 1049 -557 1061 619
rect 1003 -569 1061 -557
rect 1261 619 1319 631
rect 1261 -557 1273 619
rect 1307 -557 1319 619
rect 1261 -569 1319 -557
rect 1519 619 1577 631
rect 1519 -557 1531 619
rect 1565 -557 1577 619
rect 1519 -569 1577 -557
rect 1777 619 1835 631
rect 1777 -557 1789 619
rect 1823 -557 1835 619
rect 1777 -569 1835 -557
rect 2035 619 2093 631
rect 2035 -557 2047 619
rect 2081 -557 2093 619
rect 2035 -569 2093 -557
rect 2293 619 2351 631
rect 2293 -557 2305 619
rect 2339 -557 2351 619
rect 2293 -569 2351 -557
<< mvndiffc >>
rect -2339 -557 -2305 619
rect -2081 -557 -2047 619
rect -1823 -557 -1789 619
rect -1565 -557 -1531 619
rect -1307 -557 -1273 619
rect -1049 -557 -1015 619
rect -791 -557 -757 619
rect -533 -557 -499 619
rect -275 -557 -241 619
rect -17 -557 17 619
rect 241 -557 275 619
rect 499 -557 533 619
rect 757 -557 791 619
rect 1015 -557 1049 619
rect 1273 -557 1307 619
rect 1531 -557 1565 619
rect 1789 -557 1823 619
rect 2047 -557 2081 619
rect 2305 -557 2339 619
<< mvpsubdiff >>
rect -2485 779 2485 791
rect -2485 745 -2377 779
rect 2377 745 2485 779
rect -2485 733 2485 745
rect -2485 683 -2427 733
rect -2485 -683 -2473 683
rect -2439 -683 -2427 683
rect 2427 683 2485 733
rect -2485 -733 -2427 -683
rect 2427 -683 2439 683
rect 2473 -683 2485 683
rect 2427 -733 2485 -683
rect -2485 -745 2485 -733
rect -2485 -779 -2377 -745
rect 2377 -779 2485 -745
rect -2485 -791 2485 -779
<< mvpsubdiffcont >>
rect -2377 745 2377 779
rect -2473 -683 -2439 683
rect 2439 -683 2473 683
rect -2377 -779 2377 -745
<< poly >>
rect -2293 631 -2093 657
rect -2035 631 -1835 657
rect -1777 631 -1577 657
rect -1519 631 -1319 657
rect -1261 631 -1061 657
rect -1003 631 -803 657
rect -745 631 -545 657
rect -487 631 -287 657
rect -229 631 -29 657
rect 29 631 229 657
rect 287 631 487 657
rect 545 631 745 657
rect 803 631 1003 657
rect 1061 631 1261 657
rect 1319 631 1519 657
rect 1577 631 1777 657
rect 1835 631 2035 657
rect 2093 631 2293 657
rect -2293 -607 -2093 -569
rect -2293 -641 -2277 -607
rect -2109 -641 -2093 -607
rect -2293 -657 -2093 -641
rect -2035 -607 -1835 -569
rect -2035 -641 -2019 -607
rect -1851 -641 -1835 -607
rect -2035 -657 -1835 -641
rect -1777 -607 -1577 -569
rect -1777 -641 -1761 -607
rect -1593 -641 -1577 -607
rect -1777 -657 -1577 -641
rect -1519 -607 -1319 -569
rect -1519 -641 -1503 -607
rect -1335 -641 -1319 -607
rect -1519 -657 -1319 -641
rect -1261 -607 -1061 -569
rect -1261 -641 -1245 -607
rect -1077 -641 -1061 -607
rect -1261 -657 -1061 -641
rect -1003 -607 -803 -569
rect -1003 -641 -987 -607
rect -819 -641 -803 -607
rect -1003 -657 -803 -641
rect -745 -607 -545 -569
rect -745 -641 -729 -607
rect -561 -641 -545 -607
rect -745 -657 -545 -641
rect -487 -607 -287 -569
rect -487 -641 -471 -607
rect -303 -641 -287 -607
rect -487 -657 -287 -641
rect -229 -607 -29 -569
rect -229 -641 -213 -607
rect -45 -641 -29 -607
rect -229 -657 -29 -641
rect 29 -607 229 -569
rect 29 -641 45 -607
rect 213 -641 229 -607
rect 29 -657 229 -641
rect 287 -607 487 -569
rect 287 -641 303 -607
rect 471 -641 487 -607
rect 287 -657 487 -641
rect 545 -607 745 -569
rect 545 -641 561 -607
rect 729 -641 745 -607
rect 545 -657 745 -641
rect 803 -607 1003 -569
rect 803 -641 819 -607
rect 987 -641 1003 -607
rect 803 -657 1003 -641
rect 1061 -607 1261 -569
rect 1061 -641 1077 -607
rect 1245 -641 1261 -607
rect 1061 -657 1261 -641
rect 1319 -607 1519 -569
rect 1319 -641 1335 -607
rect 1503 -641 1519 -607
rect 1319 -657 1519 -641
rect 1577 -607 1777 -569
rect 1577 -641 1593 -607
rect 1761 -641 1777 -607
rect 1577 -657 1777 -641
rect 1835 -607 2035 -569
rect 1835 -641 1851 -607
rect 2019 -641 2035 -607
rect 1835 -657 2035 -641
rect 2093 -607 2293 -569
rect 2093 -641 2109 -607
rect 2277 -641 2293 -607
rect 2093 -657 2293 -641
<< polycont >>
rect -2277 -641 -2109 -607
rect -2019 -641 -1851 -607
rect -1761 -641 -1593 -607
rect -1503 -641 -1335 -607
rect -1245 -641 -1077 -607
rect -987 -641 -819 -607
rect -729 -641 -561 -607
rect -471 -641 -303 -607
rect -213 -641 -45 -607
rect 45 -641 213 -607
rect 303 -641 471 -607
rect 561 -641 729 -607
rect 819 -641 987 -607
rect 1077 -641 1245 -607
rect 1335 -641 1503 -607
rect 1593 -641 1761 -607
rect 1851 -641 2019 -607
rect 2109 -641 2277 -607
<< locali >>
rect -2473 745 -2377 779
rect 2377 745 2473 779
rect -2473 683 -2439 745
rect 2439 683 2473 745
rect -2339 619 -2305 635
rect -2339 -573 -2305 -557
rect -2081 619 -2047 635
rect -2081 -573 -2047 -557
rect -1823 619 -1789 635
rect -1823 -573 -1789 -557
rect -1565 619 -1531 635
rect -1565 -573 -1531 -557
rect -1307 619 -1273 635
rect -1307 -573 -1273 -557
rect -1049 619 -1015 635
rect -1049 -573 -1015 -557
rect -791 619 -757 635
rect -791 -573 -757 -557
rect -533 619 -499 635
rect -533 -573 -499 -557
rect -275 619 -241 635
rect -275 -573 -241 -557
rect -17 619 17 635
rect -17 -573 17 -557
rect 241 619 275 635
rect 241 -573 275 -557
rect 499 619 533 635
rect 499 -573 533 -557
rect 757 619 791 635
rect 757 -573 791 -557
rect 1015 619 1049 635
rect 1015 -573 1049 -557
rect 1273 619 1307 635
rect 1273 -573 1307 -557
rect 1531 619 1565 635
rect 1531 -573 1565 -557
rect 1789 619 1823 635
rect 1789 -573 1823 -557
rect 2047 619 2081 635
rect 2047 -573 2081 -557
rect 2305 619 2339 635
rect 2305 -573 2339 -557
rect -2293 -641 -2277 -607
rect -2109 -641 -2093 -607
rect -2035 -641 -2019 -607
rect -1851 -641 -1835 -607
rect -1777 -641 -1761 -607
rect -1593 -641 -1577 -607
rect -1519 -641 -1503 -607
rect -1335 -641 -1319 -607
rect -1261 -641 -1245 -607
rect -1077 -641 -1061 -607
rect -1003 -641 -987 -607
rect -819 -641 -803 -607
rect -745 -641 -729 -607
rect -561 -641 -545 -607
rect -487 -641 -471 -607
rect -303 -641 -287 -607
rect -229 -641 -213 -607
rect -45 -641 -29 -607
rect 29 -641 45 -607
rect 213 -641 229 -607
rect 287 -641 303 -607
rect 471 -641 487 -607
rect 545 -641 561 -607
rect 729 -641 745 -607
rect 803 -641 819 -607
rect 987 -641 1003 -607
rect 1061 -641 1077 -607
rect 1245 -641 1261 -607
rect 1319 -641 1335 -607
rect 1503 -641 1519 -607
rect 1577 -641 1593 -607
rect 1761 -641 1777 -607
rect 1835 -641 1851 -607
rect 2019 -641 2035 -607
rect 2093 -641 2109 -607
rect 2277 -641 2293 -607
rect -2473 -745 -2439 -683
rect 2439 -745 2473 -683
rect -2473 -779 -2377 -745
rect 2377 -779 2473 -745
<< viali >>
rect -2339 -557 -2305 619
rect -2081 -557 -2047 619
rect -1823 -557 -1789 619
rect -1565 -557 -1531 619
rect -1307 -557 -1273 619
rect -1049 -557 -1015 619
rect -791 -557 -757 619
rect -533 -557 -499 619
rect -275 -557 -241 619
rect -17 -557 17 619
rect 241 -557 275 619
rect 499 -557 533 619
rect 757 -557 791 619
rect 1015 -557 1049 619
rect 1273 -557 1307 619
rect 1531 -557 1565 619
rect 1789 -557 1823 619
rect 2047 -557 2081 619
rect 2305 -557 2339 619
rect -2277 -641 -2109 -607
rect -2019 -641 -1851 -607
rect -1761 -641 -1593 -607
rect -1503 -641 -1335 -607
rect -1245 -641 -1077 -607
rect -987 -641 -819 -607
rect -729 -641 -561 -607
rect -471 -641 -303 -607
rect -213 -641 -45 -607
rect 45 -641 213 -607
rect 303 -641 471 -607
rect 561 -641 729 -607
rect 819 -641 987 -607
rect 1077 -641 1245 -607
rect 1335 -641 1503 -607
rect 1593 -641 1761 -607
rect 1851 -641 2019 -607
rect 2109 -641 2277 -607
<< metal1 >>
rect -2345 619 -2299 631
rect -2345 -557 -2339 619
rect -2305 -557 -2299 619
rect -2345 -569 -2299 -557
rect -2087 619 -2041 631
rect -2087 -557 -2081 619
rect -2047 -557 -2041 619
rect -2087 -569 -2041 -557
rect -1829 619 -1783 631
rect -1829 -557 -1823 619
rect -1789 -557 -1783 619
rect -1829 -569 -1783 -557
rect -1571 619 -1525 631
rect -1571 -557 -1565 619
rect -1531 -557 -1525 619
rect -1571 -569 -1525 -557
rect -1313 619 -1267 631
rect -1313 -557 -1307 619
rect -1273 -557 -1267 619
rect -1313 -569 -1267 -557
rect -1055 619 -1009 631
rect -1055 -557 -1049 619
rect -1015 -557 -1009 619
rect -1055 -569 -1009 -557
rect -797 619 -751 631
rect -797 -557 -791 619
rect -757 -557 -751 619
rect -797 -569 -751 -557
rect -539 619 -493 631
rect -539 -557 -533 619
rect -499 -557 -493 619
rect -539 -569 -493 -557
rect -281 619 -235 631
rect -281 -557 -275 619
rect -241 -557 -235 619
rect -281 -569 -235 -557
rect -23 619 23 631
rect -23 -557 -17 619
rect 17 -557 23 619
rect -23 -569 23 -557
rect 235 619 281 631
rect 235 -557 241 619
rect 275 -557 281 619
rect 235 -569 281 -557
rect 493 619 539 631
rect 493 -557 499 619
rect 533 -557 539 619
rect 493 -569 539 -557
rect 751 619 797 631
rect 751 -557 757 619
rect 791 -557 797 619
rect 751 -569 797 -557
rect 1009 619 1055 631
rect 1009 -557 1015 619
rect 1049 -557 1055 619
rect 1009 -569 1055 -557
rect 1267 619 1313 631
rect 1267 -557 1273 619
rect 1307 -557 1313 619
rect 1267 -569 1313 -557
rect 1525 619 1571 631
rect 1525 -557 1531 619
rect 1565 -557 1571 619
rect 1525 -569 1571 -557
rect 1783 619 1829 631
rect 1783 -557 1789 619
rect 1823 -557 1829 619
rect 1783 -569 1829 -557
rect 2041 619 2087 631
rect 2041 -557 2047 619
rect 2081 -557 2087 619
rect 2041 -569 2087 -557
rect 2299 619 2345 631
rect 2299 -557 2305 619
rect 2339 -557 2345 619
rect 2299 -569 2345 -557
rect -2289 -607 -2097 -601
rect -2289 -641 -2277 -607
rect -2109 -641 -2097 -607
rect -2289 -647 -2097 -641
rect -2031 -607 -1839 -601
rect -2031 -641 -2019 -607
rect -1851 -641 -1839 -607
rect -2031 -647 -1839 -641
rect -1773 -607 -1581 -601
rect -1773 -641 -1761 -607
rect -1593 -641 -1581 -607
rect -1773 -647 -1581 -641
rect -1515 -607 -1323 -601
rect -1515 -641 -1503 -607
rect -1335 -641 -1323 -607
rect -1515 -647 -1323 -641
rect -1257 -607 -1065 -601
rect -1257 -641 -1245 -607
rect -1077 -641 -1065 -607
rect -1257 -647 -1065 -641
rect -999 -607 -807 -601
rect -999 -641 -987 -607
rect -819 -641 -807 -607
rect -999 -647 -807 -641
rect -741 -607 -549 -601
rect -741 -641 -729 -607
rect -561 -641 -549 -607
rect -741 -647 -549 -641
rect -483 -607 -291 -601
rect -483 -641 -471 -607
rect -303 -641 -291 -607
rect -483 -647 -291 -641
rect -225 -607 -33 -601
rect -225 -641 -213 -607
rect -45 -641 -33 -607
rect -225 -647 -33 -641
rect 33 -607 225 -601
rect 33 -641 45 -607
rect 213 -641 225 -607
rect 33 -647 225 -641
rect 291 -607 483 -601
rect 291 -641 303 -607
rect 471 -641 483 -607
rect 291 -647 483 -641
rect 549 -607 741 -601
rect 549 -641 561 -607
rect 729 -641 741 -607
rect 549 -647 741 -641
rect 807 -607 999 -601
rect 807 -641 819 -607
rect 987 -641 999 -607
rect 807 -647 999 -641
rect 1065 -607 1257 -601
rect 1065 -641 1077 -607
rect 1245 -641 1257 -607
rect 1065 -647 1257 -641
rect 1323 -607 1515 -601
rect 1323 -641 1335 -607
rect 1503 -641 1515 -607
rect 1323 -647 1515 -641
rect 1581 -607 1773 -601
rect 1581 -641 1593 -607
rect 1761 -641 1773 -607
rect 1581 -647 1773 -641
rect 1839 -607 2031 -601
rect 1839 -641 1851 -607
rect 2019 -641 2031 -607
rect 1839 -647 2031 -641
rect 2097 -607 2289 -601
rect 2097 -641 2109 -607
rect 2277 -641 2289 -607
rect 2097 -647 2289 -641
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -2456 -762 2456 762
string parameters w 6 l 1 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
