magic
tech sky130B
magscale 1 2
timestamp 1648056542
<< mvnmos >>
rect 0 0 100 200
<< mvndiff >>
rect -80 170 0 200
rect -80 30 -60 170
rect -20 30 0 170
rect -80 0 0 30
rect 100 170 180 200
rect 100 30 120 170
rect 160 30 180 170
rect 100 0 180 30
<< mvndiffc >>
rect -60 30 -20 170
rect 120 30 160 170
<< mvpsubdiff >>
rect 180 180 320 200
rect 180 20 230 180
rect 270 20 320 180
rect 180 0 320 20
<< mvpsubdiffcont >>
rect 230 20 270 180
<< poly >>
rect 0 200 100 230
rect 0 -50 100 0
rect 0 -90 20 -50
rect 80 -90 100 -50
rect 0 -110 100 -90
<< polycont >>
rect 20 -90 80 -50
<< locali >>
rect -70 175 -10 190
rect -70 25 -60 175
rect -20 25 -10 175
rect -70 10 -10 25
rect 110 170 170 190
rect 110 30 120 170
rect 160 30 170 170
rect 110 10 170 30
rect 210 180 290 190
rect 210 20 230 180
rect 270 20 290 180
rect 210 10 290 20
rect 0 -50 100 -30
rect 0 -90 20 -50
rect 80 -90 100 -50
rect 0 -110 100 -90
<< viali >>
rect -60 170 -20 175
rect -60 30 -20 170
rect -60 25 -20 30
rect 120 30 160 170
rect 230 20 270 180
rect 20 -90 80 -50
<< metal1 >>
rect -70 190 -30 230
rect -70 175 -10 190
rect -70 25 -60 175
rect -20 25 -10 175
rect 110 170 170 190
rect 110 156 120 170
rect 80 44 120 156
rect -70 10 -10 25
rect 110 30 120 44
rect 160 156 170 170
rect 220 180 280 230
rect 160 44 190 156
rect 160 30 170 44
rect 110 10 170 30
rect 220 20 230 180
rect 270 20 280 180
rect -70 -170 -30 10
rect 0 -40 100 -30
rect 0 -100 20 -40
rect 80 -100 100 -40
rect 0 -110 100 -100
rect 220 -100 280 20
rect 220 -180 280 -170
<< via1 >>
rect 20 -50 80 -40
rect 20 -90 80 -50
rect 20 -100 80 -90
rect 220 -170 280 -100
<< reram >>
rect 90 56 180 146
<< metal2 >>
rect 80 146 190 156
rect 80 130 90 146
rect -80 70 90 130
rect 80 56 90 70
rect 180 130 190 146
rect 180 70 320 130
rect 180 56 190 70
rect 80 44 190 56
rect -70 -140 -30 40
rect 0 -40 100 -30
rect 0 -100 20 -40
rect 80 -100 100 -40
rect 0 -110 100 -100
rect 210 -140 220 -100
rect -80 -170 220 -140
rect 280 -140 290 -100
rect 280 -170 320 -140
rect -70 -240 -30 -170
<< via2 >>
rect 20 -100 80 -40
<< metal3 >>
rect 0 -40 100 -30
rect 0 -50 20 -40
rect -80 -100 20 -50
rect 80 -50 100 -40
rect 80 -100 320 -50
rect -80 -110 320 -100
<< labels >>
rlabel metal2 -80 100 -80 100 7 row
port 1 w
rlabel metal1 -50 -170 -50 -170 5 col
port 2 s
rlabel metal3 -80 -80 -80 -80 7 WL
port 3 w
rlabel metal1 250 -170 250 -170 5 body
port 4 s
<< end >>
