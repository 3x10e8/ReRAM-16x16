magic
tech sky130A
magscale 1 2
timestamp 1620666330
<< pwell >>
rect -3811 -827 3811 827
<< mvnmos >>
rect -3583 -631 -3383 569
rect -3325 -631 -3125 569
rect -3067 -631 -2867 569
rect -2809 -631 -2609 569
rect -2551 -631 -2351 569
rect -2293 -631 -2093 569
rect -2035 -631 -1835 569
rect -1777 -631 -1577 569
rect -1519 -631 -1319 569
rect -1261 -631 -1061 569
rect -1003 -631 -803 569
rect -745 -631 -545 569
rect -487 -631 -287 569
rect -229 -631 -29 569
rect 29 -631 229 569
rect 287 -631 487 569
rect 545 -631 745 569
rect 803 -631 1003 569
rect 1061 -631 1261 569
rect 1319 -631 1519 569
rect 1577 -631 1777 569
rect 1835 -631 2035 569
rect 2093 -631 2293 569
rect 2351 -631 2551 569
rect 2609 -631 2809 569
rect 2867 -631 3067 569
rect 3125 -631 3325 569
rect 3383 -631 3583 569
<< mvndiff >>
rect -3641 557 -3583 569
rect -3641 -619 -3629 557
rect -3595 -619 -3583 557
rect -3641 -631 -3583 -619
rect -3383 557 -3325 569
rect -3383 -619 -3371 557
rect -3337 -619 -3325 557
rect -3383 -631 -3325 -619
rect -3125 557 -3067 569
rect -3125 -619 -3113 557
rect -3079 -619 -3067 557
rect -3125 -631 -3067 -619
rect -2867 557 -2809 569
rect -2867 -619 -2855 557
rect -2821 -619 -2809 557
rect -2867 -631 -2809 -619
rect -2609 557 -2551 569
rect -2609 -619 -2597 557
rect -2563 -619 -2551 557
rect -2609 -631 -2551 -619
rect -2351 557 -2293 569
rect -2351 -619 -2339 557
rect -2305 -619 -2293 557
rect -2351 -631 -2293 -619
rect -2093 557 -2035 569
rect -2093 -619 -2081 557
rect -2047 -619 -2035 557
rect -2093 -631 -2035 -619
rect -1835 557 -1777 569
rect -1835 -619 -1823 557
rect -1789 -619 -1777 557
rect -1835 -631 -1777 -619
rect -1577 557 -1519 569
rect -1577 -619 -1565 557
rect -1531 -619 -1519 557
rect -1577 -631 -1519 -619
rect -1319 557 -1261 569
rect -1319 -619 -1307 557
rect -1273 -619 -1261 557
rect -1319 -631 -1261 -619
rect -1061 557 -1003 569
rect -1061 -619 -1049 557
rect -1015 -619 -1003 557
rect -1061 -631 -1003 -619
rect -803 557 -745 569
rect -803 -619 -791 557
rect -757 -619 -745 557
rect -803 -631 -745 -619
rect -545 557 -487 569
rect -545 -619 -533 557
rect -499 -619 -487 557
rect -545 -631 -487 -619
rect -287 557 -229 569
rect -287 -619 -275 557
rect -241 -619 -229 557
rect -287 -631 -229 -619
rect -29 557 29 569
rect -29 -619 -17 557
rect 17 -619 29 557
rect -29 -631 29 -619
rect 229 557 287 569
rect 229 -619 241 557
rect 275 -619 287 557
rect 229 -631 287 -619
rect 487 557 545 569
rect 487 -619 499 557
rect 533 -619 545 557
rect 487 -631 545 -619
rect 745 557 803 569
rect 745 -619 757 557
rect 791 -619 803 557
rect 745 -631 803 -619
rect 1003 557 1061 569
rect 1003 -619 1015 557
rect 1049 -619 1061 557
rect 1003 -631 1061 -619
rect 1261 557 1319 569
rect 1261 -619 1273 557
rect 1307 -619 1319 557
rect 1261 -631 1319 -619
rect 1519 557 1577 569
rect 1519 -619 1531 557
rect 1565 -619 1577 557
rect 1519 -631 1577 -619
rect 1777 557 1835 569
rect 1777 -619 1789 557
rect 1823 -619 1835 557
rect 1777 -631 1835 -619
rect 2035 557 2093 569
rect 2035 -619 2047 557
rect 2081 -619 2093 557
rect 2035 -631 2093 -619
rect 2293 557 2351 569
rect 2293 -619 2305 557
rect 2339 -619 2351 557
rect 2293 -631 2351 -619
rect 2551 557 2609 569
rect 2551 -619 2563 557
rect 2597 -619 2609 557
rect 2551 -631 2609 -619
rect 2809 557 2867 569
rect 2809 -619 2821 557
rect 2855 -619 2867 557
rect 2809 -631 2867 -619
rect 3067 557 3125 569
rect 3067 -619 3079 557
rect 3113 -619 3125 557
rect 3067 -631 3125 -619
rect 3325 557 3383 569
rect 3325 -619 3337 557
rect 3371 -619 3383 557
rect 3325 -631 3383 -619
rect 3583 557 3641 569
rect 3583 -619 3595 557
rect 3629 -619 3641 557
rect 3583 -631 3641 -619
<< mvndiffc >>
rect -3629 -619 -3595 557
rect -3371 -619 -3337 557
rect -3113 -619 -3079 557
rect -2855 -619 -2821 557
rect -2597 -619 -2563 557
rect -2339 -619 -2305 557
rect -2081 -619 -2047 557
rect -1823 -619 -1789 557
rect -1565 -619 -1531 557
rect -1307 -619 -1273 557
rect -1049 -619 -1015 557
rect -791 -619 -757 557
rect -533 -619 -499 557
rect -275 -619 -241 557
rect -17 -619 17 557
rect 241 -619 275 557
rect 499 -619 533 557
rect 757 -619 791 557
rect 1015 -619 1049 557
rect 1273 -619 1307 557
rect 1531 -619 1565 557
rect 1789 -619 1823 557
rect 2047 -619 2081 557
rect 2305 -619 2339 557
rect 2563 -619 2597 557
rect 2821 -619 2855 557
rect 3079 -619 3113 557
rect 3337 -619 3371 557
rect 3595 -619 3629 557
<< mvpsubdiff >>
rect -3775 779 3775 791
rect -3775 745 -3667 779
rect 3667 745 3775 779
rect -3775 733 3775 745
rect -3775 683 -3717 733
rect -3775 -683 -3763 683
rect -3729 -683 -3717 683
rect 3717 683 3775 733
rect -3775 -733 -3717 -683
rect 3717 -683 3729 683
rect 3763 -683 3775 683
rect 3717 -733 3775 -683
rect -3775 -745 3775 -733
rect -3775 -779 -3667 -745
rect 3667 -779 3775 -745
rect -3775 -791 3775 -779
<< mvpsubdiffcont >>
rect -3667 745 3667 779
rect -3763 -683 -3729 683
rect 3729 -683 3763 683
rect -3667 -779 3667 -745
<< poly >>
rect -3583 641 -3383 657
rect -3583 607 -3567 641
rect -3399 607 -3383 641
rect -3583 569 -3383 607
rect -3325 641 -3125 657
rect -3325 607 -3309 641
rect -3141 607 -3125 641
rect -3325 569 -3125 607
rect -3067 641 -2867 657
rect -3067 607 -3051 641
rect -2883 607 -2867 641
rect -3067 569 -2867 607
rect -2809 641 -2609 657
rect -2809 607 -2793 641
rect -2625 607 -2609 641
rect -2809 569 -2609 607
rect -2551 641 -2351 657
rect -2551 607 -2535 641
rect -2367 607 -2351 641
rect -2551 569 -2351 607
rect -2293 641 -2093 657
rect -2293 607 -2277 641
rect -2109 607 -2093 641
rect -2293 569 -2093 607
rect -2035 641 -1835 657
rect -2035 607 -2019 641
rect -1851 607 -1835 641
rect -2035 569 -1835 607
rect -1777 641 -1577 657
rect -1777 607 -1761 641
rect -1593 607 -1577 641
rect -1777 569 -1577 607
rect -1519 641 -1319 657
rect -1519 607 -1503 641
rect -1335 607 -1319 641
rect -1519 569 -1319 607
rect -1261 641 -1061 657
rect -1261 607 -1245 641
rect -1077 607 -1061 641
rect -1261 569 -1061 607
rect -1003 641 -803 657
rect -1003 607 -987 641
rect -819 607 -803 641
rect -1003 569 -803 607
rect -745 641 -545 657
rect -745 607 -729 641
rect -561 607 -545 641
rect -745 569 -545 607
rect -487 641 -287 657
rect -487 607 -471 641
rect -303 607 -287 641
rect -487 569 -287 607
rect -229 641 -29 657
rect -229 607 -213 641
rect -45 607 -29 641
rect -229 569 -29 607
rect 29 641 229 657
rect 29 607 45 641
rect 213 607 229 641
rect 29 569 229 607
rect 287 641 487 657
rect 287 607 303 641
rect 471 607 487 641
rect 287 569 487 607
rect 545 641 745 657
rect 545 607 561 641
rect 729 607 745 641
rect 545 569 745 607
rect 803 641 1003 657
rect 803 607 819 641
rect 987 607 1003 641
rect 803 569 1003 607
rect 1061 641 1261 657
rect 1061 607 1077 641
rect 1245 607 1261 641
rect 1061 569 1261 607
rect 1319 641 1519 657
rect 1319 607 1335 641
rect 1503 607 1519 641
rect 1319 569 1519 607
rect 1577 641 1777 657
rect 1577 607 1593 641
rect 1761 607 1777 641
rect 1577 569 1777 607
rect 1835 641 2035 657
rect 1835 607 1851 641
rect 2019 607 2035 641
rect 1835 569 2035 607
rect 2093 641 2293 657
rect 2093 607 2109 641
rect 2277 607 2293 641
rect 2093 569 2293 607
rect 2351 641 2551 657
rect 2351 607 2367 641
rect 2535 607 2551 641
rect 2351 569 2551 607
rect 2609 641 2809 657
rect 2609 607 2625 641
rect 2793 607 2809 641
rect 2609 569 2809 607
rect 2867 641 3067 657
rect 2867 607 2883 641
rect 3051 607 3067 641
rect 2867 569 3067 607
rect 3125 641 3325 657
rect 3125 607 3141 641
rect 3309 607 3325 641
rect 3125 569 3325 607
rect 3383 641 3583 657
rect 3383 607 3399 641
rect 3567 607 3583 641
rect 3383 569 3583 607
rect -3583 -657 -3383 -631
rect -3325 -657 -3125 -631
rect -3067 -657 -2867 -631
rect -2809 -657 -2609 -631
rect -2551 -657 -2351 -631
rect -2293 -657 -2093 -631
rect -2035 -657 -1835 -631
rect -1777 -657 -1577 -631
rect -1519 -657 -1319 -631
rect -1261 -657 -1061 -631
rect -1003 -657 -803 -631
rect -745 -657 -545 -631
rect -487 -657 -287 -631
rect -229 -657 -29 -631
rect 29 -657 229 -631
rect 287 -657 487 -631
rect 545 -657 745 -631
rect 803 -657 1003 -631
rect 1061 -657 1261 -631
rect 1319 -657 1519 -631
rect 1577 -657 1777 -631
rect 1835 -657 2035 -631
rect 2093 -657 2293 -631
rect 2351 -657 2551 -631
rect 2609 -657 2809 -631
rect 2867 -657 3067 -631
rect 3125 -657 3325 -631
rect 3383 -657 3583 -631
<< polycont >>
rect -3567 607 -3399 641
rect -3309 607 -3141 641
rect -3051 607 -2883 641
rect -2793 607 -2625 641
rect -2535 607 -2367 641
rect -2277 607 -2109 641
rect -2019 607 -1851 641
rect -1761 607 -1593 641
rect -1503 607 -1335 641
rect -1245 607 -1077 641
rect -987 607 -819 641
rect -729 607 -561 641
rect -471 607 -303 641
rect -213 607 -45 641
rect 45 607 213 641
rect 303 607 471 641
rect 561 607 729 641
rect 819 607 987 641
rect 1077 607 1245 641
rect 1335 607 1503 641
rect 1593 607 1761 641
rect 1851 607 2019 641
rect 2109 607 2277 641
rect 2367 607 2535 641
rect 2625 607 2793 641
rect 2883 607 3051 641
rect 3141 607 3309 641
rect 3399 607 3567 641
<< locali >>
rect -3763 745 -3667 779
rect 3667 745 3763 779
rect -3763 683 -3729 745
rect 3729 683 3763 745
rect -3583 607 -3567 641
rect -3399 607 -3383 641
rect -3325 607 -3309 641
rect -3141 607 -3125 641
rect -3067 607 -3051 641
rect -2883 607 -2867 641
rect -2809 607 -2793 641
rect -2625 607 -2609 641
rect -2551 607 -2535 641
rect -2367 607 -2351 641
rect -2293 607 -2277 641
rect -2109 607 -2093 641
rect -2035 607 -2019 641
rect -1851 607 -1835 641
rect -1777 607 -1761 641
rect -1593 607 -1577 641
rect -1519 607 -1503 641
rect -1335 607 -1319 641
rect -1261 607 -1245 641
rect -1077 607 -1061 641
rect -1003 607 -987 641
rect -819 607 -803 641
rect -745 607 -729 641
rect -561 607 -545 641
rect -487 607 -471 641
rect -303 607 -287 641
rect -229 607 -213 641
rect -45 607 -29 641
rect 29 607 45 641
rect 213 607 229 641
rect 287 607 303 641
rect 471 607 487 641
rect 545 607 561 641
rect 729 607 745 641
rect 803 607 819 641
rect 987 607 1003 641
rect 1061 607 1077 641
rect 1245 607 1261 641
rect 1319 607 1335 641
rect 1503 607 1519 641
rect 1577 607 1593 641
rect 1761 607 1777 641
rect 1835 607 1851 641
rect 2019 607 2035 641
rect 2093 607 2109 641
rect 2277 607 2293 641
rect 2351 607 2367 641
rect 2535 607 2551 641
rect 2609 607 2625 641
rect 2793 607 2809 641
rect 2867 607 2883 641
rect 3051 607 3067 641
rect 3125 607 3141 641
rect 3309 607 3325 641
rect 3383 607 3399 641
rect 3567 607 3583 641
rect -3629 557 -3595 573
rect -3629 -635 -3595 -619
rect -3371 557 -3337 573
rect -3371 -635 -3337 -619
rect -3113 557 -3079 573
rect -3113 -635 -3079 -619
rect -2855 557 -2821 573
rect -2855 -635 -2821 -619
rect -2597 557 -2563 573
rect -2597 -635 -2563 -619
rect -2339 557 -2305 573
rect -2339 -635 -2305 -619
rect -2081 557 -2047 573
rect -2081 -635 -2047 -619
rect -1823 557 -1789 573
rect -1823 -635 -1789 -619
rect -1565 557 -1531 573
rect -1565 -635 -1531 -619
rect -1307 557 -1273 573
rect -1307 -635 -1273 -619
rect -1049 557 -1015 573
rect -1049 -635 -1015 -619
rect -791 557 -757 573
rect -791 -635 -757 -619
rect -533 557 -499 573
rect -533 -635 -499 -619
rect -275 557 -241 573
rect -275 -635 -241 -619
rect -17 557 17 573
rect -17 -635 17 -619
rect 241 557 275 573
rect 241 -635 275 -619
rect 499 557 533 573
rect 499 -635 533 -619
rect 757 557 791 573
rect 757 -635 791 -619
rect 1015 557 1049 573
rect 1015 -635 1049 -619
rect 1273 557 1307 573
rect 1273 -635 1307 -619
rect 1531 557 1565 573
rect 1531 -635 1565 -619
rect 1789 557 1823 573
rect 1789 -635 1823 -619
rect 2047 557 2081 573
rect 2047 -635 2081 -619
rect 2305 557 2339 573
rect 2305 -635 2339 -619
rect 2563 557 2597 573
rect 2563 -635 2597 -619
rect 2821 557 2855 573
rect 2821 -635 2855 -619
rect 3079 557 3113 573
rect 3079 -635 3113 -619
rect 3337 557 3371 573
rect 3337 -635 3371 -619
rect 3595 557 3629 573
rect 3595 -635 3629 -619
rect -3763 -745 -3729 -683
rect 3729 -745 3763 -683
rect -3763 -779 -3667 -745
rect 3667 -779 3763 -745
<< viali >>
rect -3567 607 -3399 641
rect -3309 607 -3141 641
rect -3051 607 -2883 641
rect -2793 607 -2625 641
rect -2535 607 -2367 641
rect -2277 607 -2109 641
rect -2019 607 -1851 641
rect -1761 607 -1593 641
rect -1503 607 -1335 641
rect -1245 607 -1077 641
rect -987 607 -819 641
rect -729 607 -561 641
rect -471 607 -303 641
rect -213 607 -45 641
rect 45 607 213 641
rect 303 607 471 641
rect 561 607 729 641
rect 819 607 987 641
rect 1077 607 1245 641
rect 1335 607 1503 641
rect 1593 607 1761 641
rect 1851 607 2019 641
rect 2109 607 2277 641
rect 2367 607 2535 641
rect 2625 607 2793 641
rect 2883 607 3051 641
rect 3141 607 3309 641
rect 3399 607 3567 641
rect -3629 -619 -3595 557
rect -3371 -619 -3337 557
rect -3113 -619 -3079 557
rect -2855 -619 -2821 557
rect -2597 -619 -2563 557
rect -2339 -619 -2305 557
rect -2081 -619 -2047 557
rect -1823 -619 -1789 557
rect -1565 -619 -1531 557
rect -1307 -619 -1273 557
rect -1049 -619 -1015 557
rect -791 -619 -757 557
rect -533 -619 -499 557
rect -275 -619 -241 557
rect -17 -619 17 557
rect 241 -619 275 557
rect 499 -619 533 557
rect 757 -619 791 557
rect 1015 -619 1049 557
rect 1273 -619 1307 557
rect 1531 -619 1565 557
rect 1789 -619 1823 557
rect 2047 -619 2081 557
rect 2305 -619 2339 557
rect 2563 -619 2597 557
rect 2821 -619 2855 557
rect 3079 -619 3113 557
rect 3337 -619 3371 557
rect 3595 -619 3629 557
<< metal1 >>
rect -3579 641 -3387 647
rect -3579 607 -3567 641
rect -3399 607 -3387 641
rect -3579 601 -3387 607
rect -3321 641 -3129 647
rect -3321 607 -3309 641
rect -3141 607 -3129 641
rect -3321 601 -3129 607
rect -3063 641 -2871 647
rect -3063 607 -3051 641
rect -2883 607 -2871 641
rect -3063 601 -2871 607
rect -2805 641 -2613 647
rect -2805 607 -2793 641
rect -2625 607 -2613 641
rect -2805 601 -2613 607
rect -2547 641 -2355 647
rect -2547 607 -2535 641
rect -2367 607 -2355 641
rect -2547 601 -2355 607
rect -2289 641 -2097 647
rect -2289 607 -2277 641
rect -2109 607 -2097 641
rect -2289 601 -2097 607
rect -2031 641 -1839 647
rect -2031 607 -2019 641
rect -1851 607 -1839 641
rect -2031 601 -1839 607
rect -1773 641 -1581 647
rect -1773 607 -1761 641
rect -1593 607 -1581 641
rect -1773 601 -1581 607
rect -1515 641 -1323 647
rect -1515 607 -1503 641
rect -1335 607 -1323 641
rect -1515 601 -1323 607
rect -1257 641 -1065 647
rect -1257 607 -1245 641
rect -1077 607 -1065 641
rect -1257 601 -1065 607
rect -999 641 -807 647
rect -999 607 -987 641
rect -819 607 -807 641
rect -999 601 -807 607
rect -741 641 -549 647
rect -741 607 -729 641
rect -561 607 -549 641
rect -741 601 -549 607
rect -483 641 -291 647
rect -483 607 -471 641
rect -303 607 -291 641
rect -483 601 -291 607
rect -225 641 -33 647
rect -225 607 -213 641
rect -45 607 -33 641
rect -225 601 -33 607
rect 33 641 225 647
rect 33 607 45 641
rect 213 607 225 641
rect 33 601 225 607
rect 291 641 483 647
rect 291 607 303 641
rect 471 607 483 641
rect 291 601 483 607
rect 549 641 741 647
rect 549 607 561 641
rect 729 607 741 641
rect 549 601 741 607
rect 807 641 999 647
rect 807 607 819 641
rect 987 607 999 641
rect 807 601 999 607
rect 1065 641 1257 647
rect 1065 607 1077 641
rect 1245 607 1257 641
rect 1065 601 1257 607
rect 1323 641 1515 647
rect 1323 607 1335 641
rect 1503 607 1515 641
rect 1323 601 1515 607
rect 1581 641 1773 647
rect 1581 607 1593 641
rect 1761 607 1773 641
rect 1581 601 1773 607
rect 1839 641 2031 647
rect 1839 607 1851 641
rect 2019 607 2031 641
rect 1839 601 2031 607
rect 2097 641 2289 647
rect 2097 607 2109 641
rect 2277 607 2289 641
rect 2097 601 2289 607
rect 2355 641 2547 647
rect 2355 607 2367 641
rect 2535 607 2547 641
rect 2355 601 2547 607
rect 2613 641 2805 647
rect 2613 607 2625 641
rect 2793 607 2805 641
rect 2613 601 2805 607
rect 2871 641 3063 647
rect 2871 607 2883 641
rect 3051 607 3063 641
rect 2871 601 3063 607
rect 3129 641 3321 647
rect 3129 607 3141 641
rect 3309 607 3321 641
rect 3129 601 3321 607
rect 3387 641 3579 647
rect 3387 607 3399 641
rect 3567 607 3579 641
rect 3387 601 3579 607
rect -3635 557 -3589 569
rect -3635 -619 -3629 557
rect -3595 -619 -3589 557
rect -3635 -631 -3589 -619
rect -3377 557 -3331 569
rect -3377 -619 -3371 557
rect -3337 -619 -3331 557
rect -3377 -631 -3331 -619
rect -3119 557 -3073 569
rect -3119 -619 -3113 557
rect -3079 -619 -3073 557
rect -3119 -631 -3073 -619
rect -2861 557 -2815 569
rect -2861 -619 -2855 557
rect -2821 -619 -2815 557
rect -2861 -631 -2815 -619
rect -2603 557 -2557 569
rect -2603 -619 -2597 557
rect -2563 -619 -2557 557
rect -2603 -631 -2557 -619
rect -2345 557 -2299 569
rect -2345 -619 -2339 557
rect -2305 -619 -2299 557
rect -2345 -631 -2299 -619
rect -2087 557 -2041 569
rect -2087 -619 -2081 557
rect -2047 -619 -2041 557
rect -2087 -631 -2041 -619
rect -1829 557 -1783 569
rect -1829 -619 -1823 557
rect -1789 -619 -1783 557
rect -1829 -631 -1783 -619
rect -1571 557 -1525 569
rect -1571 -619 -1565 557
rect -1531 -619 -1525 557
rect -1571 -631 -1525 -619
rect -1313 557 -1267 569
rect -1313 -619 -1307 557
rect -1273 -619 -1267 557
rect -1313 -631 -1267 -619
rect -1055 557 -1009 569
rect -1055 -619 -1049 557
rect -1015 -619 -1009 557
rect -1055 -631 -1009 -619
rect -797 557 -751 569
rect -797 -619 -791 557
rect -757 -619 -751 557
rect -797 -631 -751 -619
rect -539 557 -493 569
rect -539 -619 -533 557
rect -499 -619 -493 557
rect -539 -631 -493 -619
rect -281 557 -235 569
rect -281 -619 -275 557
rect -241 -619 -235 557
rect -281 -631 -235 -619
rect -23 557 23 569
rect -23 -619 -17 557
rect 17 -619 23 557
rect -23 -631 23 -619
rect 235 557 281 569
rect 235 -619 241 557
rect 275 -619 281 557
rect 235 -631 281 -619
rect 493 557 539 569
rect 493 -619 499 557
rect 533 -619 539 557
rect 493 -631 539 -619
rect 751 557 797 569
rect 751 -619 757 557
rect 791 -619 797 557
rect 751 -631 797 -619
rect 1009 557 1055 569
rect 1009 -619 1015 557
rect 1049 -619 1055 557
rect 1009 -631 1055 -619
rect 1267 557 1313 569
rect 1267 -619 1273 557
rect 1307 -619 1313 557
rect 1267 -631 1313 -619
rect 1525 557 1571 569
rect 1525 -619 1531 557
rect 1565 -619 1571 557
rect 1525 -631 1571 -619
rect 1783 557 1829 569
rect 1783 -619 1789 557
rect 1823 -619 1829 557
rect 1783 -631 1829 -619
rect 2041 557 2087 569
rect 2041 -619 2047 557
rect 2081 -619 2087 557
rect 2041 -631 2087 -619
rect 2299 557 2345 569
rect 2299 -619 2305 557
rect 2339 -619 2345 557
rect 2299 -631 2345 -619
rect 2557 557 2603 569
rect 2557 -619 2563 557
rect 2597 -619 2603 557
rect 2557 -631 2603 -619
rect 2815 557 2861 569
rect 2815 -619 2821 557
rect 2855 -619 2861 557
rect 2815 -631 2861 -619
rect 3073 557 3119 569
rect 3073 -619 3079 557
rect 3113 -619 3119 557
rect 3073 -631 3119 -619
rect 3331 557 3377 569
rect 3331 -619 3337 557
rect 3371 -619 3377 557
rect 3331 -631 3377 -619
rect 3589 557 3635 569
rect 3589 -619 3595 557
rect 3629 -619 3635 557
rect 3589 -631 3635 -619
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -3746 -762 3746 762
string parameters w 6 l 1 m 1 nf 28 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
