magic
tech sky130B
timestamp 1647920407
<< nwell >>
rect -30 -2124 1110 -1924
<< mvnmos >>
rect 1190 -2059 1240 -1959
rect 1285 -2059 1335 -1959
rect 1380 -2059 1430 -1959
rect 1475 -2059 1525 -1959
rect 1570 -2059 1620 -1959
rect 1780 -2059 1830 -1959
rect 1875 -2059 1925 -1959
rect 1970 -2059 2020 -1959
rect 2065 -2059 2115 -1959
rect 2160 -2059 2210 -1959
rect 2255 -2059 2305 -1959
rect 2350 -2059 2400 -1959
<< mvpmos >>
rect 55 -2059 105 -1959
rect 150 -2059 200 -1959
rect 245 -2059 295 -1959
rect 340 -2059 390 -1959
rect 435 -2059 485 -1959
rect 530 -2059 580 -1959
rect 625 -2059 675 -1959
rect 720 -2059 770 -1959
rect 815 -2059 865 -1959
rect 910 -2059 960 -1959
<< mvndiff >>
rect 1145 -1985 1190 -1959
rect 1145 -2044 1155 -1985
rect 1180 -2044 1190 -1985
rect 1145 -2059 1190 -2044
rect 1240 -1974 1285 -1959
rect 1240 -2044 1250 -1974
rect 1275 -2044 1285 -1974
rect 1240 -2059 1285 -2044
rect 1335 -1985 1380 -1959
rect 1335 -2044 1345 -1985
rect 1370 -2044 1380 -1985
rect 1335 -2059 1380 -2044
rect 1430 -1974 1475 -1959
rect 1430 -2044 1440 -1974
rect 1465 -2044 1475 -1974
rect 1430 -2059 1475 -2044
rect 1525 -1983 1570 -1959
rect 1525 -2044 1535 -1983
rect 1560 -2044 1570 -1983
rect 1525 -2059 1570 -2044
rect 1620 -1979 1665 -1959
rect 1620 -2044 1630 -1979
rect 1655 -2044 1665 -1979
rect 1735 -1979 1780 -1959
rect 1735 -2044 1745 -1979
rect 1770 -2044 1780 -1979
rect 1620 -2059 1665 -2044
rect 1735 -2059 1780 -2044
rect 1830 -1974 1875 -1959
rect 1830 -2044 1840 -1974
rect 1865 -2044 1875 -1974
rect 1830 -2059 1875 -2044
rect 1925 -1986 1970 -1959
rect 1925 -2044 1935 -1986
rect 1960 -2044 1970 -1986
rect 1925 -2059 1970 -2044
rect 2020 -1974 2065 -1959
rect 2020 -2044 2030 -1974
rect 2055 -2044 2065 -1974
rect 2020 -2059 2065 -2044
rect 2115 -1984 2160 -1959
rect 2115 -2044 2125 -1984
rect 2150 -2044 2160 -1984
rect 2115 -2059 2160 -2044
rect 2210 -1974 2255 -1959
rect 2210 -2044 2220 -1974
rect 2245 -2044 2255 -1974
rect 2210 -2059 2255 -2044
rect 2305 -1984 2350 -1959
rect 2305 -2044 2315 -1984
rect 2340 -2044 2350 -1984
rect 2305 -2059 2350 -2044
rect 2400 -1974 2445 -1959
rect 2400 -2044 2410 -1974
rect 2435 -2044 2445 -1974
rect 2400 -2059 2445 -2044
<< mvpdiff >>
rect 10 -1979 55 -1959
rect 10 -2044 20 -1979
rect 45 -2044 55 -1979
rect 10 -2059 55 -2044
rect 105 -1974 150 -1959
rect 105 -2044 115 -1974
rect 140 -2044 150 -1974
rect 105 -2059 150 -2044
rect 200 -1986 245 -1959
rect 200 -2044 210 -1986
rect 235 -2044 245 -1986
rect 200 -2059 245 -2044
rect 295 -1974 340 -1959
rect 295 -2044 305 -1974
rect 330 -2044 340 -1974
rect 295 -2059 340 -2044
rect 390 -1985 435 -1959
rect 390 -2044 400 -1985
rect 425 -2044 435 -1985
rect 390 -2059 435 -2044
rect 485 -1974 530 -1959
rect 485 -2044 495 -1974
rect 520 -2044 530 -1974
rect 485 -2059 530 -2044
rect 580 -1985 625 -1959
rect 580 -2044 590 -1985
rect 615 -2044 625 -1985
rect 580 -2059 625 -2044
rect 675 -1974 720 -1959
rect 675 -2044 685 -1974
rect 710 -2044 720 -1974
rect 675 -2059 720 -2044
rect 770 -1988 815 -1959
rect 770 -2044 780 -1988
rect 805 -2044 815 -1988
rect 770 -2059 815 -2044
rect 865 -1974 910 -1959
rect 865 -2044 875 -1974
rect 900 -2044 910 -1974
rect 865 -2059 910 -2044
rect 960 -1979 1005 -1959
rect 960 -2044 970 -1979
rect 995 -2044 1005 -1979
rect 960 -2059 1005 -2044
<< mvndiffc >>
rect 1155 -2044 1180 -1985
rect 1250 -2044 1275 -1974
rect 1345 -2044 1370 -1985
rect 1440 -2044 1465 -1974
rect 1535 -2044 1560 -1983
rect 1630 -2044 1655 -1979
rect 1745 -2044 1770 -1979
rect 1840 -2044 1865 -1974
rect 1935 -2044 1960 -1986
rect 2030 -2044 2055 -1974
rect 2125 -2044 2150 -1984
rect 2220 -2044 2245 -1974
rect 2315 -2044 2340 -1984
rect 2410 -2044 2435 -1974
<< mvpdiffc >>
rect 20 -2044 45 -1979
rect 115 -2044 140 -1974
rect 210 -2044 235 -1986
rect 305 -2044 330 -1974
rect 400 -2044 425 -1985
rect 495 -2044 520 -1974
rect 590 -2044 615 -1985
rect 685 -2044 710 -1974
rect 780 -2044 805 -1988
rect 875 -2044 900 -1974
rect 970 -2044 995 -1979
<< mvpsubdiff >>
rect 1665 -1986 1735 -1959
rect 1665 -2044 1681 -1986
rect 1719 -2044 1735 -1986
rect 1665 -2059 1735 -2044
<< mvnsubdiff >>
rect 1005 -1974 1075 -1959
rect 1005 -2044 1030 -1974
rect 1060 -2044 1075 -1974
rect 1005 -2059 1075 -2044
<< mvpsubdiffcont >>
rect 1681 -2044 1719 -1986
<< mvnsubdiffcont >>
rect 1030 -2044 1060 -1974
<< poly >>
rect 55 -1959 105 -1944
rect 150 -1959 200 -1944
rect 245 -1959 295 -1944
rect 340 -1959 390 -1944
rect 435 -1959 485 -1944
rect 530 -1959 580 -1944
rect 625 -1959 675 -1944
rect 720 -1959 770 -1944
rect 815 -1959 865 -1944
rect 910 -1959 960 -1944
rect 1190 -1959 1240 -1944
rect 1285 -1959 1335 -1944
rect 1380 -1959 1430 -1944
rect 1475 -1959 1525 -1944
rect 1570 -1959 1620 -1944
rect 1780 -1959 1830 -1944
rect 1875 -1959 1925 -1944
rect 1970 -1959 2020 -1944
rect 2065 -1959 2115 -1944
rect 2160 -1959 2210 -1944
rect 2255 -1959 2305 -1944
rect 2350 -1959 2400 -1944
rect 55 -2084 105 -2059
rect 55 -2114 65 -2084
rect 95 -2114 105 -2084
rect 55 -2119 105 -2114
rect 150 -2084 200 -2059
rect 150 -2114 160 -2084
rect 190 -2114 200 -2084
rect 150 -2119 200 -2114
rect 245 -2084 295 -2059
rect 245 -2114 255 -2084
rect 285 -2114 295 -2084
rect 245 -2119 295 -2114
rect 340 -2084 390 -2059
rect 340 -2114 350 -2084
rect 380 -2114 390 -2084
rect 340 -2119 390 -2114
rect 435 -2084 485 -2059
rect 435 -2114 445 -2084
rect 475 -2114 485 -2084
rect 435 -2119 485 -2114
rect 530 -2084 580 -2059
rect 530 -2114 540 -2084
rect 570 -2114 580 -2084
rect 530 -2119 580 -2114
rect 625 -2084 675 -2059
rect 625 -2114 635 -2084
rect 665 -2114 675 -2084
rect 625 -2119 675 -2114
rect 720 -2084 770 -2059
rect 720 -2114 730 -2084
rect 760 -2114 770 -2084
rect 720 -2119 770 -2114
rect 815 -2084 865 -2059
rect 815 -2114 825 -2084
rect 855 -2114 865 -2084
rect 815 -2119 865 -2114
rect 910 -2084 960 -2059
rect 910 -2114 920 -2084
rect 950 -2114 960 -2084
rect 910 -2119 960 -2114
rect 1190 -2084 1240 -2059
rect 1190 -2114 1200 -2084
rect 1230 -2114 1240 -2084
rect 1190 -2119 1240 -2114
rect 1285 -2084 1335 -2059
rect 1285 -2114 1295 -2084
rect 1325 -2114 1335 -2084
rect 1285 -2119 1335 -2114
rect 1380 -2084 1430 -2059
rect 1380 -2114 1390 -2084
rect 1420 -2114 1430 -2084
rect 1380 -2119 1430 -2114
rect 1475 -2084 1525 -2059
rect 1475 -2114 1485 -2084
rect 1515 -2114 1525 -2084
rect 1475 -2119 1525 -2114
rect 1570 -2084 1620 -2059
rect 1570 -2114 1580 -2084
rect 1610 -2114 1620 -2084
rect 1570 -2119 1620 -2114
rect 1780 -2084 1830 -2059
rect 1780 -2114 1790 -2084
rect 1820 -2114 1830 -2084
rect 1780 -2119 1830 -2114
rect 1875 -2084 1925 -2059
rect 1875 -2114 1885 -2084
rect 1915 -2114 1925 -2084
rect 1875 -2119 1925 -2114
rect 1970 -2084 2020 -2059
rect 1970 -2114 1980 -2084
rect 2010 -2114 2020 -2084
rect 1970 -2119 2020 -2114
rect 2065 -2084 2115 -2059
rect 2065 -2114 2075 -2084
rect 2105 -2114 2115 -2084
rect 2065 -2119 2115 -2114
rect 2160 -2084 2210 -2059
rect 2160 -2114 2170 -2084
rect 2200 -2114 2210 -2084
rect 2160 -2119 2210 -2114
rect 2255 -2084 2305 -2059
rect 2255 -2114 2265 -2084
rect 2295 -2114 2305 -2084
rect 2255 -2119 2305 -2114
rect 2350 -2084 2400 -2059
rect 2350 -2114 2360 -2084
rect 2390 -2114 2400 -2084
rect 2350 -2119 2400 -2114
<< polycont >>
rect 65 -2114 95 -2084
rect 160 -2114 190 -2084
rect 255 -2114 285 -2084
rect 350 -2114 380 -2084
rect 445 -2114 475 -2084
rect 540 -2114 570 -2084
rect 635 -2114 665 -2084
rect 730 -2114 760 -2084
rect 825 -2114 855 -2084
rect 920 -2114 950 -2084
rect 1200 -2114 1230 -2084
rect 1295 -2114 1325 -2084
rect 1390 -2114 1420 -2084
rect 1485 -2114 1515 -2084
rect 1580 -2114 1610 -2084
rect 1790 -2114 1820 -2084
rect 1885 -2114 1915 -2084
rect 1980 -2114 2010 -2084
rect 2075 -2114 2105 -2084
rect 2170 -2114 2200 -2084
rect 2265 -2114 2295 -2084
rect 2360 -2114 2390 -2084
<< locali >>
rect 68 -1958 905 -1941
rect 1145 -1958 1660 -1941
rect 15 -1979 50 -1969
rect 15 -2044 20 -1979
rect 45 -2044 50 -1979
rect 15 -2054 50 -2044
rect 110 -1974 145 -1958
rect 110 -2044 115 -1974
rect 140 -2044 145 -1974
rect 300 -1974 335 -1958
rect 110 -2054 145 -2044
rect 205 -1979 240 -1975
rect 205 -2044 210 -1979
rect 235 -2044 240 -1979
rect 205 -2054 240 -2044
rect 300 -2044 305 -1974
rect 330 -2044 335 -1974
rect 490 -1974 525 -1958
rect 300 -2054 335 -2044
rect 395 -1979 430 -1975
rect 395 -2044 400 -1979
rect 425 -2044 430 -1979
rect 395 -2054 430 -2044
rect 490 -2044 495 -1974
rect 520 -2044 525 -1974
rect 680 -1974 715 -1958
rect 490 -2054 525 -2044
rect 585 -1979 620 -1975
rect 585 -2044 590 -1979
rect 615 -2044 620 -1979
rect 585 -2054 620 -2044
rect 680 -2044 685 -1974
rect 710 -2044 715 -1974
rect 870 -1974 905 -1958
rect 680 -2054 715 -2044
rect 775 -1979 810 -1975
rect 775 -2044 780 -1979
rect 805 -2044 810 -1979
rect 775 -2054 810 -2044
rect 870 -2044 875 -1974
rect 900 -2044 905 -1974
rect 870 -2054 905 -2044
rect 965 -1979 1000 -1969
rect 965 -2044 970 -1979
rect 995 -2044 1000 -1979
rect 965 -2054 1000 -2044
rect 1020 -1974 1070 -1964
rect 1020 -2044 1030 -1974
rect 1060 -2044 1070 -1974
rect 1245 -1974 1280 -1958
rect 1020 -2054 1070 -2044
rect 1150 -1979 1185 -1975
rect 1150 -2044 1155 -1979
rect 1180 -2044 1185 -1979
rect 1150 -2054 1185 -2044
rect 1245 -2044 1250 -1974
rect 1275 -2044 1280 -1974
rect 1435 -1974 1470 -1958
rect 1245 -2054 1280 -2044
rect 1340 -1979 1375 -1975
rect 1340 -2044 1345 -1979
rect 1370 -2044 1375 -1979
rect 1340 -2054 1375 -2044
rect 1435 -2044 1440 -1974
rect 1465 -2044 1470 -1974
rect 1435 -2054 1470 -2044
rect 1530 -2044 1535 -1975
rect 1560 -2044 1565 -1975
rect 1530 -2054 1565 -2044
rect 1625 -1979 1660 -1958
rect 1835 -1958 2440 -1941
rect 1625 -2044 1630 -1979
rect 1655 -2044 1660 -1979
rect 1625 -2054 1660 -2044
rect 1677 -2044 1681 -1975
rect 1719 -2044 1723 -1975
rect 1677 -2054 1723 -2044
rect 1740 -1979 1775 -1964
rect 1740 -2044 1745 -1979
rect 1770 -2044 1775 -1979
rect 1740 -2054 1775 -2044
rect 1835 -1974 1870 -1958
rect 1835 -2044 1840 -1974
rect 1865 -2044 1870 -1974
rect 2025 -1974 2060 -1958
rect 1835 -2054 1870 -2044
rect 1930 -1979 1965 -1975
rect 1930 -2044 1935 -1979
rect 1960 -2044 1965 -1979
rect 1930 -2054 1965 -2044
rect 2025 -2044 2030 -1974
rect 2055 -2044 2060 -1974
rect 2215 -1974 2250 -1958
rect 2025 -2054 2060 -2044
rect 2120 -1979 2155 -1975
rect 2120 -2044 2125 -1979
rect 2150 -2044 2155 -1979
rect 2120 -2054 2155 -2044
rect 2215 -2044 2220 -1974
rect 2245 -2044 2250 -1974
rect 2405 -1974 2440 -1958
rect 2215 -2054 2250 -2044
rect 2310 -1979 2345 -1975
rect 2310 -2044 2315 -1979
rect 2340 -2044 2345 -1979
rect 2310 -2054 2345 -2044
rect 2405 -2044 2410 -1974
rect 2435 -2044 2440 -1974
rect 2405 -2054 2440 -2044
rect 60 -2084 100 -2074
rect 60 -2114 65 -2084
rect 95 -2114 100 -2084
rect 60 -2124 100 -2114
rect 155 -2084 195 -2074
rect 155 -2114 160 -2084
rect 190 -2114 195 -2084
rect 155 -2124 195 -2114
rect 250 -2084 290 -2074
rect 250 -2114 255 -2084
rect 285 -2114 290 -2084
rect 250 -2124 290 -2114
rect 345 -2084 385 -2074
rect 345 -2114 350 -2084
rect 380 -2114 385 -2084
rect 345 -2124 385 -2114
rect 440 -2084 480 -2074
rect 440 -2114 445 -2084
rect 475 -2114 480 -2084
rect 440 -2124 480 -2114
rect 535 -2084 575 -2074
rect 630 -2084 670 -2074
rect 725 -2084 765 -2074
rect 820 -2084 860 -2074
rect 915 -2084 955 -2074
rect 535 -2114 540 -2084
rect 570 -2114 635 -2084
rect 665 -2114 730 -2084
rect 760 -2114 825 -2084
rect 855 -2114 920 -2084
rect 950 -2114 955 -2084
rect 535 -2124 575 -2114
rect 630 -2124 670 -2114
rect 725 -2124 765 -2114
rect 820 -2124 860 -2114
rect 915 -2124 955 -2114
rect 1195 -2084 1235 -2074
rect 1195 -2114 1200 -2084
rect 1230 -2114 1235 -2084
rect 1195 -2124 1235 -2114
rect 1290 -2084 1330 -2074
rect 1290 -2114 1295 -2084
rect 1325 -2114 1330 -2084
rect 1290 -2124 1330 -2114
rect 1385 -2084 1425 -2074
rect 1385 -2114 1390 -2084
rect 1420 -2114 1425 -2084
rect 1385 -2124 1425 -2114
rect 1480 -2084 1520 -2074
rect 1575 -2084 1615 -2074
rect 1480 -2114 1485 -2084
rect 1515 -2114 1580 -2084
rect 1610 -2114 1615 -2084
rect 1480 -2124 1520 -2114
rect 1575 -2124 1615 -2114
rect 1785 -2084 1825 -2074
rect 1785 -2114 1790 -2084
rect 1820 -2114 1825 -2084
rect 1785 -2124 1825 -2114
rect 1880 -2084 1920 -2074
rect 1880 -2114 1885 -2084
rect 1915 -2114 1920 -2084
rect 1880 -2124 1920 -2114
rect 1975 -2084 2015 -2074
rect 1975 -2114 1980 -2084
rect 2010 -2114 2015 -2084
rect 1975 -2124 2015 -2114
rect 2070 -2084 2110 -2074
rect 2165 -2084 2205 -2074
rect 2070 -2114 2075 -2084
rect 2105 -2114 2170 -2084
rect 2200 -2114 2205 -2084
rect 2070 -2124 2110 -2114
rect 2165 -2124 2205 -2114
rect 2260 -2084 2300 -2074
rect 2355 -2084 2395 -2074
rect 2260 -2114 2265 -2084
rect 2295 -2114 2360 -2084
rect 2390 -2114 2395 -2084
rect 2260 -2124 2300 -2114
rect 2355 -2124 2395 -2114
<< viali >>
rect 20 -2044 45 -1979
rect 210 -1986 235 -1979
rect 210 -2044 235 -1986
rect 400 -1985 425 -1979
rect 400 -2044 425 -1985
rect 590 -1985 615 -1979
rect 590 -2044 615 -1985
rect 780 -1988 805 -1979
rect 780 -2044 805 -1988
rect 970 -2044 995 -1979
rect 1030 -2044 1060 -1974
rect 1155 -1985 1180 -1979
rect 1155 -2044 1180 -1985
rect 1345 -1985 1370 -1979
rect 1345 -2044 1370 -1985
rect 1535 -1983 1560 -1975
rect 1535 -2044 1560 -1983
rect 1681 -1986 1719 -1975
rect 1681 -2044 1719 -1986
rect 1745 -2044 1770 -1979
rect 1935 -1986 1960 -1979
rect 1935 -2044 1960 -1986
rect 2125 -1984 2150 -1979
rect 2125 -2044 2150 -1984
rect 2315 -1984 2340 -1979
rect 2315 -2044 2340 -1984
rect 65 -2114 95 -2084
rect 160 -2114 190 -2084
rect 255 -2114 285 -2084
rect 350 -2114 380 -2084
rect 445 -2114 475 -2084
rect 540 -2114 570 -2084
rect 635 -2114 665 -2084
rect 730 -2114 760 -2084
rect 825 -2114 855 -2084
rect 920 -2114 950 -2084
rect 1200 -2114 1230 -2084
rect 1295 -2114 1325 -2084
rect 1390 -2114 1420 -2084
rect 1485 -2114 1515 -2084
rect 1580 -2114 1610 -2084
rect 1790 -2114 1820 -2084
rect 1885 -2114 1915 -2084
rect 1980 -2114 2010 -2084
rect 2075 -2114 2105 -2084
rect 2170 -2114 2200 -2084
rect 2265 -2114 2295 -2084
rect 2360 -2114 2390 -2084
<< metal1 >>
rect 15 -1979 50 -1969
rect 15 -2054 50 -2044
rect 205 -1979 240 -1969
rect 205 -2054 240 -2044
rect 395 -1979 430 -1969
rect 395 -2054 430 -2044
rect 540 -2074 570 -1924
rect 590 -1939 615 -1924
rect 780 -1939 805 -1924
rect 970 -1939 995 -1924
rect 590 -1954 995 -1939
rect 590 -1969 615 -1954
rect 780 -1969 805 -1954
rect 970 -1969 995 -1954
rect 585 -1979 620 -1969
rect 585 -2044 590 -1979
rect 615 -2044 620 -1979
rect 585 -2054 620 -2044
rect 775 -1979 810 -1969
rect 775 -2044 780 -1979
rect 805 -2044 810 -1979
rect 775 -2054 810 -2044
rect 965 -1979 1000 -1969
rect 965 -2044 970 -1979
rect 995 -2044 1000 -1979
rect 965 -2054 1000 -2044
rect 1025 -1974 1065 -1924
rect 1025 -2044 1030 -1974
rect 1060 -2044 1065 -1974
rect 60 -2084 100 -2074
rect 60 -2114 65 -2084
rect 95 -2114 100 -2084
rect 60 -2124 100 -2114
rect 155 -2084 195 -2074
rect 155 -2114 160 -2084
rect 190 -2114 195 -2084
rect 155 -2124 195 -2114
rect 250 -2084 290 -2074
rect 250 -2114 255 -2084
rect 285 -2114 290 -2084
rect 250 -2124 290 -2114
rect 345 -2084 385 -2074
rect 345 -2114 350 -2084
rect 380 -2114 385 -2084
rect 345 -2124 385 -2114
rect 440 -2084 480 -2074
rect 440 -2114 445 -2084
rect 475 -2114 480 -2084
rect 440 -2124 480 -2114
rect 535 -2084 575 -2074
rect 535 -2114 540 -2084
rect 570 -2114 575 -2084
rect 535 -2124 575 -2114
rect 590 -2124 615 -2054
rect 630 -2084 670 -2074
rect 630 -2114 635 -2084
rect 665 -2114 670 -2084
rect 630 -2124 670 -2114
rect 725 -2084 765 -2074
rect 725 -2114 730 -2084
rect 760 -2114 765 -2084
rect 725 -2124 765 -2114
rect 780 -2124 805 -2054
rect 820 -2084 860 -2074
rect 820 -2114 825 -2084
rect 855 -2114 860 -2084
rect 820 -2124 860 -2114
rect 915 -2084 955 -2074
rect 915 -2114 920 -2084
rect 950 -2114 955 -2084
rect 915 -2124 955 -2114
rect 970 -2124 995 -2054
rect 1025 -2124 1065 -2044
rect 1150 -1979 1185 -1969
rect 1150 -2054 1185 -2044
rect 1340 -1979 1375 -1969
rect 1340 -2054 1375 -2044
rect 1485 -2074 1515 -1924
rect 1535 -1939 1560 -1924
rect 1530 -1975 1565 -1939
rect 1530 -2044 1535 -1975
rect 1560 -2044 1565 -1975
rect 1530 -2054 1565 -2044
rect 1195 -2084 1235 -2074
rect 1195 -2114 1200 -2084
rect 1230 -2114 1235 -2084
rect 1195 -2124 1235 -2114
rect 1290 -2084 1330 -2074
rect 1290 -2114 1295 -2084
rect 1325 -2114 1330 -2084
rect 1290 -2124 1330 -2114
rect 1385 -2084 1425 -2074
rect 1385 -2114 1390 -2084
rect 1420 -2114 1425 -2084
rect 1385 -2124 1425 -2114
rect 1480 -2084 1520 -2074
rect 1480 -2114 1485 -2084
rect 1515 -2114 1520 -2084
rect 1480 -2124 1520 -2114
rect 1535 -2124 1560 -2054
rect 1580 -2074 1610 -1924
rect 1677 -1975 1723 -1924
rect 2125 -1969 2150 -1924
rect 1677 -2044 1681 -1975
rect 1719 -2044 1723 -1975
rect 1575 -2084 1615 -2074
rect 1575 -2114 1580 -2084
rect 1610 -2114 1615 -2084
rect 1575 -2124 1615 -2114
rect 1677 -2124 1723 -2044
rect 1740 -1979 1775 -1969
rect 1740 -2054 1775 -2044
rect 1930 -1979 1965 -1969
rect 1930 -2054 1965 -2044
rect 2120 -1979 2155 -1969
rect 2120 -2044 2125 -1979
rect 2150 -2044 2155 -1979
rect 2120 -2054 2155 -2044
rect 1785 -2084 1825 -2074
rect 1785 -2114 1790 -2084
rect 1820 -2114 1825 -2084
rect 1785 -2124 1825 -2114
rect 1880 -2084 1920 -2074
rect 1880 -2114 1885 -2084
rect 1915 -2114 1920 -2084
rect 1880 -2124 1920 -2114
rect 1975 -2084 2015 -2074
rect 1975 -2114 1980 -2084
rect 2010 -2114 2015 -2084
rect 1975 -2124 2015 -2114
rect 2070 -2084 2110 -2074
rect 2070 -2114 2075 -2084
rect 2105 -2114 2110 -2084
rect 2070 -2124 2110 -2114
rect 2125 -2124 2150 -2054
rect 2175 -2074 2195 -1924
rect 2315 -1969 2340 -1924
rect 2310 -1979 2345 -1969
rect 2310 -2044 2315 -1979
rect 2340 -2044 2345 -1979
rect 2310 -2054 2345 -2044
rect 2165 -2084 2205 -2074
rect 2165 -2114 2170 -2084
rect 2200 -2114 2205 -2084
rect 2165 -2124 2205 -2114
rect 2260 -2084 2300 -2074
rect 2260 -2114 2265 -2084
rect 2295 -2114 2300 -2084
rect 2260 -2124 2300 -2114
rect 2315 -2124 2340 -2054
rect 2365 -2074 2385 -1924
rect 2355 -2084 2395 -2074
rect 2355 -2114 2360 -2084
rect 2390 -2114 2395 -2084
rect 2355 -2124 2395 -2114
<< via1 >>
rect 15 -2044 20 -1979
rect 20 -2044 45 -1979
rect 45 -2044 50 -1979
rect 205 -2044 210 -1979
rect 210 -2044 235 -1979
rect 235 -2044 240 -1979
rect 395 -2044 400 -1979
rect 400 -2044 425 -1979
rect 425 -2044 430 -1979
rect 65 -2114 95 -2084
rect 160 -2114 190 -2084
rect 255 -2114 285 -2084
rect 350 -2114 380 -2084
rect 445 -2114 475 -2084
rect 1150 -2044 1155 -1979
rect 1155 -2044 1180 -1979
rect 1180 -2044 1185 -1979
rect 1340 -2044 1345 -1979
rect 1345 -2044 1370 -1979
rect 1370 -2044 1375 -1979
rect 1200 -2114 1230 -2084
rect 1295 -2114 1325 -2084
rect 1390 -2114 1420 -2084
rect 1740 -2044 1745 -1979
rect 1745 -2044 1770 -1979
rect 1770 -2044 1775 -1979
rect 1930 -2044 1935 -1979
rect 1935 -2044 1960 -1979
rect 1960 -2044 1965 -1979
rect 1790 -2114 1820 -2084
rect 1885 -2114 1915 -2084
rect 1980 -2114 2010 -2084
<< metal2 >>
rect 15 -1959 1965 -1939
rect 15 -1979 50 -1959
rect -66 -2019 15 -1999
rect 15 -2054 50 -2044
rect 205 -1979 240 -1959
rect 205 -2054 240 -2044
rect 395 -1979 430 -1959
rect 395 -2054 430 -2044
rect 1150 -1979 1185 -1959
rect 1150 -2054 1185 -2044
rect 1340 -1979 1375 -1959
rect 1340 -2054 1375 -2044
rect 1740 -1979 1775 -1959
rect 1740 -2054 1775 -2044
rect 1930 -1979 1965 -1959
rect 1930 -2054 1965 -2044
rect 60 -2084 100 -2074
rect 60 -2114 65 -2084
rect 95 -2114 100 -2084
rect 60 -2124 100 -2114
rect 155 -2084 195 -2074
rect 155 -2114 160 -2084
rect 190 -2114 195 -2084
rect 155 -2124 195 -2114
rect 250 -2084 290 -2074
rect 250 -2114 255 -2084
rect 285 -2114 290 -2084
rect 250 -2124 290 -2114
rect 345 -2084 385 -2074
rect 345 -2114 350 -2084
rect 380 -2114 385 -2084
rect 345 -2124 385 -2114
rect 440 -2084 480 -2074
rect 440 -2114 445 -2084
rect 475 -2114 480 -2084
rect 440 -2124 480 -2114
rect 1195 -2084 1235 -2074
rect 1195 -2114 1200 -2084
rect 1230 -2114 1235 -2084
rect 1195 -2124 1235 -2114
rect 1290 -2084 1330 -2074
rect 1290 -2114 1295 -2084
rect 1325 -2114 1330 -2084
rect 1290 -2124 1330 -2114
rect 1385 -2084 1425 -2074
rect 1385 -2114 1390 -2084
rect 1420 -2114 1425 -2084
rect 1385 -2124 1425 -2114
rect 1785 -2084 1825 -2074
rect 1785 -2114 1790 -2084
rect 1820 -2089 1825 -2084
rect 1880 -2084 1920 -2074
rect 1880 -2089 1885 -2084
rect 1820 -2109 1885 -2089
rect 1820 -2114 1825 -2109
rect 1785 -2124 1825 -2114
rect 1880 -2114 1885 -2109
rect 1915 -2089 1920 -2084
rect 1975 -2084 2015 -2074
rect 1975 -2089 1980 -2084
rect 1915 -2109 1980 -2089
rect 1915 -2114 1920 -2109
rect 1880 -2124 1920 -2114
rect 1975 -2114 1980 -2109
rect 2010 -2089 2015 -2084
rect 2010 -2109 2445 -2089
rect 2010 -2114 2015 -2109
rect 1975 -2124 2015 -2114
<< via2 >>
rect 65 -2114 95 -2084
rect 160 -2114 190 -2084
rect 255 -2114 285 -2084
rect 350 -2114 380 -2084
rect 445 -2114 475 -2084
rect 1200 -2114 1230 -2084
rect 1295 -2114 1325 -2084
rect 1390 -2114 1420 -2084
<< metal3 >>
rect 55 -2083 105 -2074
rect 55 -2115 64 -2083
rect 96 -2115 105 -2083
rect 55 -2124 105 -2115
rect 150 -2083 200 -2074
rect 150 -2115 159 -2083
rect 191 -2115 200 -2083
rect 150 -2124 200 -2115
rect 245 -2083 295 -2074
rect 245 -2115 254 -2083
rect 286 -2115 295 -2083
rect 245 -2124 295 -2115
rect 340 -2083 390 -2074
rect 340 -2115 349 -2083
rect 381 -2115 390 -2083
rect 340 -2124 390 -2115
rect 435 -2083 485 -2074
rect 435 -2115 444 -2083
rect 476 -2115 485 -2083
rect 435 -2124 485 -2115
rect 1190 -2084 1240 -2074
rect 1285 -2084 1335 -2074
rect 1380 -2084 1430 -2074
rect 1190 -2114 1200 -2084
rect 1230 -2114 1295 -2084
rect 1325 -2114 1390 -2084
rect 1420 -2114 2445 -2084
rect 1190 -2125 1240 -2114
rect 1285 -2125 1335 -2114
rect 1380 -2125 1430 -2114
<< via3 >>
rect 64 -2084 96 -2083
rect 64 -2114 65 -2084
rect 65 -2114 95 -2084
rect 95 -2114 96 -2084
rect 64 -2115 96 -2114
rect 159 -2084 191 -2083
rect 159 -2114 160 -2084
rect 160 -2114 190 -2084
rect 190 -2114 191 -2084
rect 159 -2115 191 -2114
rect 254 -2084 286 -2083
rect 254 -2114 255 -2084
rect 255 -2114 285 -2084
rect 285 -2114 286 -2084
rect 254 -2115 286 -2114
rect 349 -2084 381 -2083
rect 349 -2114 350 -2084
rect 350 -2114 380 -2084
rect 380 -2114 381 -2084
rect 349 -2115 381 -2114
rect 444 -2084 476 -2083
rect 444 -2114 445 -2084
rect 445 -2114 475 -2084
rect 475 -2114 476 -2084
rect 444 -2115 476 -2114
<< metal4 >>
rect 60 -2083 100 -2074
rect 60 -2115 64 -2083
rect 96 -2084 100 -2083
rect 155 -2083 195 -2074
rect 155 -2084 159 -2083
rect 96 -2114 159 -2084
rect 96 -2115 100 -2114
rect 60 -2124 100 -2115
rect 155 -2115 159 -2114
rect 191 -2084 195 -2083
rect 250 -2083 290 -2074
rect 250 -2084 254 -2083
rect 191 -2114 254 -2084
rect 191 -2115 195 -2114
rect 155 -2124 195 -2115
rect 250 -2115 254 -2114
rect 286 -2084 290 -2083
rect 345 -2083 385 -2074
rect 345 -2084 349 -2083
rect 286 -2114 349 -2084
rect 286 -2115 290 -2114
rect 250 -2124 290 -2115
rect 345 -2115 349 -2114
rect 381 -2084 385 -2083
rect 440 -2083 480 -2074
rect 440 -2084 444 -2083
rect 381 -2114 444 -2084
rect 381 -2115 385 -2114
rect 345 -2124 385 -2115
rect 440 -2115 444 -2114
rect 476 -2084 480 -2083
rect 535 -2084 575 -2074
rect 630 -2084 670 -2074
rect 725 -2084 765 -2074
rect 820 -2084 860 -2074
rect 915 -2084 955 -2074
rect 476 -2114 2445 -2084
rect 476 -2115 480 -2114
rect 440 -2124 480 -2115
rect 535 -2124 575 -2114
rect 630 -2124 670 -2114
rect 725 -2124 765 -2114
rect 820 -2124 860 -2114
rect 915 -2124 955 -2114
<< labels >>
rlabel metal1 1045 -1924 1045 -1924 1 VP
rlabel metal1 1545 -1924 1545 -1924 1 Vr-
rlabel metal1 1700 -1924 1700 -1924 1 VN
rlabel metal1 1500 -1924 1500 -1924 1 Vgn
rlabel metal1 985 -1924 985 -1924 1 Vr+
rlabel metal1 2140 -1924 2140 -1924 1 Vref
rlabel metal1 2185 -1924 2185 -1924 1 WR
rlabel metal1 2330 -1924 2330 -1924 1 Vsample
rlabel metal1 2375 -1924 2375 -1924 1 SAMPLE
rlabel metal1 555 -1924 555 -1924 1 Vgp
rlabel metal3 2445 -2099 2445 -2099 3 SWref
rlabel metal4 2445 -2094 2445 -2094 3 SWr+
rlabel metal2 2445 -2103 2445 -2103 3 SWr-
rlabel metal2 -30 -2009 -30 -2009 7 row
<< end >>
