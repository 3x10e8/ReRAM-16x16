magic
tech sky130B
timestamp 1647920282
<< nwell >>
rect -30 -789 170 351
<< mvnmos >>
rect 5 -919 105 -869
rect 5 -1014 105 -964
rect 5 -1109 105 -1059
rect 5 -1204 105 -1154
rect 5 -1299 105 -1249
rect 5 -1509 105 -1459
rect 5 -1604 105 -1554
rect 5 -1699 105 -1649
rect 5 -1794 105 -1744
rect 5 -1889 105 -1839
<< mvpmos >>
rect 5 216 105 266
rect 5 121 105 171
rect 5 26 105 76
rect 5 -69 105 -19
rect 5 -164 105 -114
rect 5 -259 105 -209
rect 5 -354 105 -304
rect 5 -449 105 -399
rect 5 -544 105 -494
rect 5 -639 105 -589
<< mvndiff >>
rect 5 -834 105 -824
rect 5 -859 31 -834
rect 90 -859 105 -834
rect 5 -869 105 -859
rect 5 -929 105 -919
rect 5 -954 20 -929
rect 90 -954 105 -929
rect 5 -964 105 -954
rect 5 -1024 105 -1014
rect 5 -1049 31 -1024
rect 90 -1049 105 -1024
rect 5 -1059 105 -1049
rect 5 -1119 105 -1109
rect 5 -1144 20 -1119
rect 90 -1144 105 -1119
rect 5 -1154 105 -1144
rect 5 -1214 105 -1204
rect 5 -1239 29 -1214
rect 90 -1239 105 -1214
rect 5 -1249 105 -1239
rect 5 -1309 105 -1299
rect 5 -1334 25 -1309
rect 90 -1334 105 -1309
rect 5 -1344 105 -1334
rect 5 -1424 105 -1414
rect 5 -1449 25 -1424
rect 90 -1449 105 -1424
rect 5 -1459 105 -1449
rect 5 -1519 105 -1509
rect 5 -1544 20 -1519
rect 90 -1544 105 -1519
rect 5 -1554 105 -1544
rect 5 -1614 105 -1604
rect 5 -1639 32 -1614
rect 90 -1639 105 -1614
rect 5 -1649 105 -1639
rect 5 -1709 105 -1699
rect 5 -1734 20 -1709
rect 90 -1734 105 -1709
rect 5 -1744 105 -1734
rect 5 -1804 105 -1794
rect 5 -1829 30 -1804
rect 90 -1829 105 -1804
rect 5 -1839 105 -1829
rect 5 -1899 105 -1889
rect 5 -1924 20 -1899
rect 90 -1924 105 -1899
rect 5 -1934 105 -1924
<< mvpdiff >>
rect 5 301 105 311
rect 5 276 25 301
rect 90 276 105 301
rect 5 266 105 276
rect 5 206 105 216
rect 5 181 20 206
rect 90 181 105 206
rect 5 171 105 181
rect 5 111 105 121
rect 5 86 32 111
rect 90 86 105 111
rect 5 76 105 86
rect 5 16 105 26
rect 5 -9 20 16
rect 90 -9 105 16
rect 5 -19 105 -9
rect 5 -79 105 -69
rect 5 -104 31 -79
rect 90 -104 105 -79
rect 5 -114 105 -104
rect 5 -174 105 -164
rect 5 -199 20 -174
rect 90 -199 105 -174
rect 5 -209 105 -199
rect 5 -269 105 -259
rect 5 -294 31 -269
rect 90 -294 105 -269
rect 5 -304 105 -294
rect 5 -364 105 -354
rect 5 -389 20 -364
rect 90 -389 105 -364
rect 5 -399 105 -389
rect 5 -459 105 -449
rect 5 -484 34 -459
rect 90 -484 105 -459
rect 5 -494 105 -484
rect 5 -554 105 -544
rect 5 -579 20 -554
rect 90 -579 105 -554
rect 5 -589 105 -579
rect 5 -649 105 -639
rect 5 -674 25 -649
rect 90 -674 105 -649
rect 5 -684 105 -674
<< mvndiffc >>
rect 31 -859 90 -834
rect 20 -954 90 -929
rect 31 -1049 90 -1024
rect 20 -1144 90 -1119
rect 29 -1239 90 -1214
rect 25 -1334 90 -1309
rect 25 -1449 90 -1424
rect 20 -1544 90 -1519
rect 32 -1639 90 -1614
rect 20 -1734 90 -1709
rect 30 -1829 90 -1804
rect 20 -1924 90 -1899
<< mvpdiffc >>
rect 25 276 90 301
rect 20 181 90 206
rect 32 86 90 111
rect 20 -9 90 16
rect 31 -104 90 -79
rect 20 -199 90 -174
rect 31 -294 90 -269
rect 20 -389 90 -364
rect 34 -484 90 -459
rect 20 -579 90 -554
rect 25 -674 90 -649
<< mvpsubdiff >>
rect 5 -1360 105 -1344
rect 5 -1398 32 -1360
rect 90 -1398 105 -1360
rect 5 -1414 105 -1398
<< mvnsubdiff >>
rect 5 -709 105 -684
rect 5 -739 20 -709
rect 90 -739 105 -709
rect 5 -754 105 -739
<< mvpsubdiffcont >>
rect 32 -1398 90 -1360
<< mvnsubdiffcont >>
rect 20 -739 90 -709
<< poly >>
rect -10 216 5 266
rect 105 256 165 266
rect 105 226 130 256
rect 160 226 165 256
rect 105 216 165 226
rect -10 121 5 171
rect 105 161 165 171
rect 105 131 130 161
rect 160 131 165 161
rect 105 121 165 131
rect -10 26 5 76
rect 105 66 165 76
rect 105 36 130 66
rect 160 36 165 66
rect 105 26 165 36
rect -10 -69 5 -19
rect 105 -29 165 -19
rect 105 -59 130 -29
rect 160 -59 165 -29
rect 105 -69 165 -59
rect -10 -164 5 -114
rect 105 -124 165 -114
rect 105 -154 130 -124
rect 160 -154 165 -124
rect 105 -164 165 -154
rect -10 -259 5 -209
rect 105 -219 165 -209
rect 105 -249 130 -219
rect 160 -249 165 -219
rect 105 -259 165 -249
rect -10 -354 5 -304
rect 105 -314 165 -304
rect 105 -344 130 -314
rect 160 -344 165 -314
rect 105 -354 165 -344
rect -10 -449 5 -399
rect 105 -409 165 -399
rect 105 -439 130 -409
rect 160 -439 165 -409
rect 105 -449 165 -439
rect -10 -544 5 -494
rect 105 -504 165 -494
rect 105 -534 130 -504
rect 160 -534 165 -504
rect 105 -544 165 -534
rect -10 -639 5 -589
rect 105 -599 165 -589
rect 105 -629 130 -599
rect 160 -629 165 -599
rect 105 -639 165 -629
rect -10 -919 5 -869
rect 105 -879 165 -869
rect 105 -909 130 -879
rect 160 -909 165 -879
rect 105 -919 165 -909
rect -10 -1014 5 -964
rect 105 -974 165 -964
rect 105 -1004 130 -974
rect 160 -1004 165 -974
rect 105 -1014 165 -1004
rect -10 -1109 5 -1059
rect 105 -1069 165 -1059
rect 105 -1099 130 -1069
rect 160 -1099 165 -1069
rect 105 -1109 165 -1099
rect -10 -1204 5 -1154
rect 105 -1164 165 -1154
rect 105 -1194 130 -1164
rect 160 -1194 165 -1164
rect 105 -1204 165 -1194
rect -10 -1299 5 -1249
rect 105 -1259 165 -1249
rect 105 -1289 130 -1259
rect 160 -1289 165 -1259
rect 105 -1299 165 -1289
rect -10 -1509 5 -1459
rect 105 -1469 165 -1459
rect 105 -1499 130 -1469
rect 160 -1499 165 -1469
rect 105 -1509 165 -1499
rect -10 -1604 5 -1554
rect 105 -1564 165 -1554
rect 105 -1594 130 -1564
rect 160 -1594 165 -1564
rect 105 -1604 165 -1594
rect -10 -1699 5 -1649
rect 105 -1659 165 -1649
rect 105 -1689 130 -1659
rect 160 -1689 165 -1659
rect 105 -1699 165 -1689
rect -10 -1794 5 -1744
rect 105 -1754 165 -1744
rect 105 -1784 130 -1754
rect 160 -1784 165 -1754
rect 105 -1794 165 -1784
rect -10 -1889 5 -1839
rect 105 -1849 165 -1839
rect 105 -1879 130 -1849
rect 160 -1879 165 -1849
rect 105 -1889 165 -1879
<< polycont >>
rect 130 226 160 256
rect 130 131 160 161
rect 130 36 160 66
rect 130 -59 160 -29
rect 130 -154 160 -124
rect 130 -249 160 -219
rect 130 -344 160 -314
rect 130 -439 160 -409
rect 130 -534 160 -504
rect 130 -629 160 -599
rect 130 -909 160 -879
rect 130 -1004 160 -974
rect 130 -1099 160 -1069
rect 130 -1194 160 -1164
rect 130 -1289 160 -1259
rect 130 -1499 160 -1469
rect 130 -1594 160 -1564
rect 130 -1689 160 -1659
rect 130 -1784 160 -1754
rect 130 -1879 160 -1849
<< locali >>
rect 15 301 100 306
rect 15 276 25 301
rect 90 276 100 301
rect 15 271 100 276
rect 120 256 170 261
rect -13 211 4 253
rect 120 226 130 256
rect 160 226 170 256
rect 120 221 170 226
rect -13 206 100 211
rect -13 181 20 206
rect 90 181 100 206
rect -13 176 100 181
rect -13 21 4 176
rect 120 161 170 166
rect 120 131 130 161
rect 160 131 170 161
rect 120 126 170 131
rect 21 111 100 116
rect 21 86 25 111
rect 90 86 100 111
rect 21 81 100 86
rect 120 66 170 71
rect 120 36 130 66
rect 160 36 170 66
rect 120 31 170 36
rect -13 16 100 21
rect -13 -9 20 16
rect 90 -9 100 16
rect -13 -14 100 -9
rect -13 -169 4 -14
rect 120 -29 170 -24
rect 120 -59 130 -29
rect 160 -59 170 -29
rect 120 -64 170 -59
rect 21 -79 100 -74
rect 21 -104 25 -79
rect 90 -104 100 -79
rect 21 -109 100 -104
rect 120 -124 170 -119
rect 120 -154 130 -124
rect 160 -154 170 -124
rect 120 -159 170 -154
rect -13 -174 100 -169
rect -13 -199 20 -174
rect 90 -199 100 -174
rect -13 -204 100 -199
rect -13 -359 4 -204
rect 120 -219 170 -214
rect 120 -249 130 -219
rect 160 -249 170 -219
rect 120 -254 170 -249
rect 21 -269 100 -264
rect 21 -294 25 -269
rect 90 -294 100 -269
rect 21 -299 100 -294
rect 130 -309 160 -254
rect 120 -314 170 -309
rect 120 -344 130 -314
rect 160 -344 170 -314
rect 120 -349 170 -344
rect -13 -364 100 -359
rect -13 -389 20 -364
rect 90 -389 100 -364
rect -13 -394 100 -389
rect -13 -549 4 -394
rect 130 -404 160 -349
rect 120 -409 170 -404
rect 120 -439 130 -409
rect 160 -439 170 -409
rect 120 -444 170 -439
rect 21 -459 100 -454
rect 21 -484 25 -459
rect 90 -484 100 -459
rect 21 -489 100 -484
rect 130 -499 160 -444
rect 120 -504 170 -499
rect 120 -534 130 -504
rect 160 -534 170 -504
rect 120 -539 170 -534
rect -13 -554 100 -549
rect -13 -579 20 -554
rect 90 -579 100 -554
rect -13 -584 100 -579
rect 130 -594 160 -539
rect 120 -599 170 -594
rect 120 -629 130 -599
rect 160 -629 170 -599
rect 120 -634 170 -629
rect 15 -649 100 -644
rect 15 -674 25 -649
rect 90 -674 100 -649
rect 15 -679 100 -674
rect 10 -709 100 -699
rect 10 -739 20 -709
rect 90 -739 100 -709
rect 10 -749 100 -739
rect -13 -924 4 -824
rect 21 -834 100 -829
rect 21 -859 25 -834
rect 90 -859 100 -834
rect 21 -864 100 -859
rect 120 -879 170 -874
rect 120 -909 130 -879
rect 160 -909 170 -879
rect 120 -914 170 -909
rect -13 -929 100 -924
rect -13 -954 20 -929
rect 90 -954 100 -929
rect -13 -959 100 -954
rect -13 -1114 4 -959
rect 120 -974 170 -969
rect 120 -1004 130 -974
rect 160 -1004 170 -974
rect 120 -1009 170 -1004
rect 21 -1024 100 -1019
rect 21 -1049 25 -1024
rect 90 -1049 100 -1024
rect 21 -1054 100 -1049
rect 120 -1069 170 -1064
rect 120 -1099 130 -1069
rect 160 -1099 170 -1069
rect 120 -1104 170 -1099
rect -13 -1119 100 -1114
rect -13 -1144 20 -1119
rect 90 -1144 100 -1119
rect -13 -1149 100 -1144
rect -13 -1304 4 -1149
rect 120 -1164 170 -1159
rect 120 -1194 130 -1164
rect 160 -1194 170 -1164
rect 120 -1199 170 -1194
rect 21 -1214 100 -1209
rect 90 -1239 100 -1214
rect 21 -1244 100 -1239
rect 130 -1254 160 -1199
rect 120 -1259 170 -1254
rect 120 -1289 130 -1259
rect 160 -1289 170 -1259
rect 120 -1294 170 -1289
rect -13 -1309 100 -1304
rect -13 -1334 25 -1309
rect 90 -1334 100 -1309
rect -13 -1339 100 -1334
rect 21 -1360 100 -1356
rect 90 -1398 100 -1360
rect 21 -1402 100 -1398
rect 10 -1424 100 -1419
rect 10 -1449 25 -1424
rect 90 -1449 100 -1424
rect 10 -1454 100 -1449
rect 120 -1469 170 -1464
rect 120 -1499 130 -1469
rect 160 -1499 170 -1469
rect 120 -1504 170 -1499
rect -13 -1519 100 -1514
rect -13 -1544 20 -1519
rect 90 -1544 100 -1519
rect -13 -1549 100 -1544
rect -13 -1704 4 -1549
rect 120 -1564 170 -1559
rect 120 -1594 130 -1564
rect 160 -1594 170 -1564
rect 120 -1599 170 -1594
rect 21 -1614 100 -1609
rect 21 -1639 25 -1614
rect 90 -1639 100 -1614
rect 21 -1644 100 -1639
rect 120 -1659 170 -1654
rect 120 -1689 130 -1659
rect 160 -1689 170 -1659
rect 120 -1694 170 -1689
rect -13 -1709 100 -1704
rect -13 -1734 20 -1709
rect 90 -1734 100 -1709
rect -13 -1739 100 -1734
rect -13 -1894 4 -1739
rect 120 -1754 170 -1749
rect 120 -1784 130 -1754
rect 160 -1784 170 -1754
rect 120 -1789 170 -1784
rect 21 -1804 100 -1799
rect 21 -1829 25 -1804
rect 90 -1829 100 -1804
rect 21 -1834 100 -1829
rect 120 -1849 170 -1844
rect 120 -1879 130 -1849
rect 160 -1879 170 -1849
rect 120 -1884 170 -1879
rect -13 -1899 100 -1894
rect -13 -1924 20 -1899
rect 90 -1924 100 -1899
rect -13 -1929 100 -1924
<< viali >>
rect 25 276 90 301
rect 130 226 160 256
rect 130 131 160 161
rect 25 86 32 111
rect 32 86 90 111
rect 130 36 160 66
rect 130 -59 160 -29
rect 25 -104 31 -79
rect 31 -104 90 -79
rect 130 -154 160 -124
rect 130 -249 160 -219
rect 25 -294 31 -269
rect 31 -294 90 -269
rect 130 -344 160 -314
rect 130 -439 160 -409
rect 25 -484 34 -459
rect 34 -484 90 -459
rect 130 -534 160 -504
rect 130 -629 160 -599
rect 25 -674 90 -649
rect 20 -739 90 -709
rect 25 -859 31 -834
rect 31 -859 90 -834
rect 130 -909 160 -879
rect 130 -1004 160 -974
rect 25 -1049 31 -1024
rect 31 -1049 90 -1024
rect 130 -1099 160 -1069
rect 130 -1194 160 -1164
rect 21 -1239 29 -1214
rect 29 -1239 90 -1214
rect 130 -1289 160 -1259
rect 21 -1398 32 -1360
rect 32 -1398 90 -1360
rect 25 -1449 90 -1424
rect 130 -1499 160 -1469
rect 20 -1544 90 -1519
rect 130 -1594 160 -1564
rect 25 -1639 32 -1614
rect 32 -1639 90 -1614
rect 130 -1689 160 -1659
rect 20 -1734 90 -1709
rect 130 -1784 160 -1754
rect 25 -1829 30 -1804
rect 30 -1829 90 -1804
rect 130 -1879 160 -1849
rect 20 -1924 90 -1899
<< metal1 >>
rect -25 351 66 371
rect 46 306 66 351
rect 15 271 25 306
rect 90 271 100 306
rect 120 256 170 261
rect 120 226 130 256
rect 160 226 170 256
rect 120 221 170 226
rect 120 161 170 166
rect 120 131 130 161
rect 160 131 170 161
rect 120 126 170 131
rect 15 81 25 116
rect 90 81 100 116
rect 120 66 170 71
rect 120 36 130 66
rect 160 36 170 66
rect 120 31 170 36
rect 120 -29 170 -24
rect 120 -59 130 -29
rect 160 -59 170 -29
rect 120 -64 170 -59
rect 15 -109 25 -74
rect 90 -109 100 -74
rect 120 -124 170 -119
rect 120 -154 130 -124
rect 160 -154 170 -124
rect 120 -159 170 -154
rect 120 -219 170 -214
rect -30 -249 130 -219
rect 160 -249 170 -219
rect 120 -254 170 -249
rect 15 -269 100 -264
rect -30 -294 25 -269
rect 90 -294 170 -269
rect -15 -459 0 -294
rect 15 -299 100 -294
rect 120 -314 170 -309
rect 120 -344 130 -314
rect 160 -344 170 -314
rect 120 -349 170 -344
rect 120 -409 170 -404
rect 120 -439 130 -409
rect 160 -439 170 -409
rect 120 -444 170 -439
rect 15 -459 100 -454
rect -30 -484 25 -459
rect 90 -484 170 -459
rect -15 -649 0 -484
rect 15 -489 100 -484
rect 120 -504 170 -499
rect 120 -534 130 -504
rect 160 -534 170 -504
rect 120 -539 170 -534
rect 120 -599 170 -594
rect 120 -629 130 -599
rect 160 -629 170 -599
rect 120 -634 170 -629
rect 15 -649 100 -644
rect -30 -674 25 -649
rect 90 -674 170 -649
rect 15 -679 100 -674
rect -30 -709 170 -704
rect -30 -739 20 -709
rect 90 -739 170 -709
rect -30 -744 170 -739
rect 15 -864 25 -829
rect 90 -864 100 -829
rect 120 -879 170 -874
rect 120 -909 130 -879
rect 160 -909 170 -879
rect 120 -914 170 -909
rect 120 -974 170 -969
rect 120 -1004 130 -974
rect 160 -1004 170 -974
rect 120 -1009 170 -1004
rect 15 -1054 25 -1019
rect 90 -1054 100 -1019
rect 120 -1069 170 -1064
rect 120 -1099 130 -1069
rect 160 -1099 170 -1069
rect 120 -1104 170 -1099
rect 120 -1164 170 -1159
rect -30 -1194 130 -1164
rect 160 -1194 170 -1164
rect 120 -1199 170 -1194
rect -15 -1214 100 -1209
rect -30 -1239 21 -1214
rect 90 -1239 170 -1214
rect -15 -1244 100 -1239
rect 120 -1259 170 -1254
rect -30 -1289 130 -1259
rect 160 -1289 170 -1259
rect 120 -1294 170 -1289
rect -30 -1360 170 -1356
rect -30 -1398 21 -1360
rect 90 -1398 170 -1360
rect -30 -1402 170 -1398
rect 15 -1454 25 -1419
rect 90 -1454 100 -1419
rect 120 -1469 170 -1464
rect 120 -1499 130 -1469
rect 160 -1499 170 -1469
rect 120 -1504 170 -1499
rect 6 -1519 100 -1513
rect -30 -1544 20 -1519
rect 90 -1544 170 -1519
rect 6 -1549 100 -1544
rect 120 -1564 170 -1559
rect 120 -1594 130 -1564
rect 160 -1594 170 -1564
rect 120 -1599 170 -1594
rect 15 -1644 25 -1609
rect 90 -1644 100 -1609
rect 120 -1659 170 -1654
rect 120 -1689 130 -1659
rect 160 -1689 170 -1659
rect 120 -1694 170 -1689
rect 6 -1709 100 -1703
rect -30 -1734 20 -1709
rect 90 -1734 170 -1709
rect 6 -1739 100 -1734
rect 120 -1754 170 -1749
rect 120 -1784 130 -1754
rect 160 -1784 170 -1754
rect 120 -1789 170 -1784
rect 15 -1834 25 -1799
rect 90 -1834 100 -1799
rect 120 -1849 170 -1844
rect 120 -1879 130 -1849
rect 160 -1879 170 -1849
rect 120 -1884 170 -1879
rect 6 -1899 100 -1893
rect -30 -1924 20 -1899
rect 90 -1924 170 -1899
rect 6 -1929 100 -1924
<< via1 >>
rect 25 301 90 306
rect 25 276 90 301
rect 25 271 90 276
rect 130 226 160 256
rect 130 131 160 161
rect 25 111 90 116
rect 25 86 90 111
rect 25 81 90 86
rect 130 36 160 66
rect 130 -59 160 -29
rect 25 -79 90 -74
rect 25 -104 90 -79
rect 25 -109 90 -104
rect 130 -154 160 -124
rect 25 -834 90 -829
rect 25 -859 90 -834
rect 25 -864 90 -859
rect 130 -909 160 -879
rect 130 -1004 160 -974
rect 25 -1024 90 -1019
rect 25 -1049 90 -1024
rect 25 -1054 90 -1049
rect 130 -1099 160 -1069
rect 25 -1424 90 -1419
rect 25 -1449 90 -1424
rect 25 -1454 90 -1449
rect 130 -1499 160 -1469
rect 130 -1594 160 -1564
rect 25 -1614 90 -1609
rect 25 -1639 90 -1614
rect 25 -1644 90 -1639
rect 130 -1689 160 -1659
rect 130 -1784 160 -1754
rect 25 -1804 90 -1799
rect 25 -1829 90 -1804
rect 25 -1834 90 -1829
rect 130 -1879 160 -1849
<< metal2 >>
rect -15 271 25 306
rect 90 271 100 306
rect -15 116 5 271
rect 120 256 170 261
rect 120 226 130 256
rect 160 226 170 256
rect 120 221 170 226
rect 120 161 170 166
rect 120 131 130 161
rect 160 131 170 161
rect 120 126 170 131
rect -15 81 25 116
rect 90 81 100 116
rect -15 -74 5 81
rect 120 66 170 71
rect 120 36 130 66
rect 160 36 170 66
rect 120 31 170 36
rect 120 -29 170 -24
rect 120 -59 130 -29
rect 160 -59 170 -29
rect 120 -64 170 -59
rect -15 -109 25 -74
rect 90 -109 100 -74
rect -15 -829 5 -109
rect 120 -124 170 -119
rect 120 -154 130 -124
rect 160 -154 170 -124
rect 120 -159 170 -154
rect -15 -864 25 -829
rect 90 -864 100 -829
rect -15 -1019 5 -864
rect 120 -879 170 -874
rect 120 -909 130 -879
rect 160 -909 170 -879
rect 120 -914 170 -909
rect 120 -974 170 -969
rect 120 -1004 130 -974
rect 160 -1004 170 -974
rect 120 -1009 170 -1004
rect -15 -1054 25 -1019
rect 90 -1054 100 -1019
rect -15 -1419 5 -1054
rect 120 -1069 170 -1064
rect 120 -1099 130 -1069
rect 160 -1099 170 -1069
rect 120 -1104 170 -1099
rect -15 -1454 25 -1419
rect 90 -1454 100 -1419
rect -15 -1609 5 -1454
rect 120 -1469 170 -1464
rect 120 -1499 130 -1469
rect 160 -1499 170 -1469
rect 120 -1504 170 -1499
rect 135 -1559 155 -1504
rect 120 -1564 170 -1559
rect 120 -1594 130 -1564
rect 160 -1594 170 -1564
rect 120 -1599 170 -1594
rect -15 -1644 25 -1609
rect 90 -1644 100 -1609
rect -15 -1799 5 -1644
rect 135 -1654 155 -1599
rect 120 -1659 170 -1654
rect 120 -1689 130 -1659
rect 160 -1689 170 -1659
rect 120 -1694 170 -1689
rect 135 -1749 155 -1694
rect 120 -1754 170 -1749
rect 120 -1784 130 -1754
rect 160 -1784 170 -1754
rect 120 -1789 170 -1784
rect -15 -1834 25 -1799
rect 90 -1834 100 -1799
rect 135 -1844 155 -1789
rect 120 -1849 170 -1844
rect 120 -1879 130 -1849
rect 160 -1879 170 -1849
rect 120 -1884 170 -1879
rect -15 -1929 5 -1893
rect 135 -1934 155 -1884
<< via2 >>
rect 130 226 160 256
rect 130 131 160 161
rect 130 36 160 66
rect 130 -59 160 -29
rect 130 -154 160 -124
rect 130 -909 160 -879
rect 130 -1004 160 -974
rect 130 -1099 160 -1069
<< metal3 >>
rect 120 257 170 266
rect 120 225 129 257
rect 161 225 170 257
rect 120 216 170 225
rect 120 162 170 171
rect 120 130 129 162
rect 161 130 170 162
rect 120 121 170 130
rect 120 67 170 76
rect 120 35 129 67
rect 161 35 170 67
rect 120 26 170 35
rect 120 -28 170 -19
rect 120 -60 129 -28
rect 161 -60 170 -28
rect 120 -69 170 -60
rect 120 -123 170 -114
rect 120 -155 129 -123
rect 161 -155 170 -123
rect 120 -164 170 -155
rect 120 -879 170 -869
rect 120 -909 130 -879
rect 160 -909 170 -879
rect 120 -919 170 -909
rect 130 -964 160 -919
rect 120 -974 170 -964
rect 120 -1004 130 -974
rect 160 -1004 170 -974
rect 120 -1014 170 -1004
rect 130 -1059 160 -1014
rect 120 -1069 170 -1059
rect 120 -1099 130 -1069
rect 160 -1099 170 -1069
rect 120 -1109 170 -1099
rect 130 -1934 160 -1109
<< via3 >>
rect 129 256 161 257
rect 129 226 130 256
rect 130 226 160 256
rect 160 226 161 256
rect 129 225 161 226
rect 129 161 161 162
rect 129 131 130 161
rect 130 131 160 161
rect 160 131 161 161
rect 129 130 161 131
rect 129 66 161 67
rect 129 36 130 66
rect 130 36 160 66
rect 160 36 161 66
rect 129 35 161 36
rect 129 -29 161 -28
rect 129 -59 130 -29
rect 130 -59 160 -29
rect 160 -59 161 -29
rect 129 -60 161 -59
rect 129 -124 161 -123
rect 129 -154 130 -124
rect 130 -154 160 -124
rect 160 -154 161 -124
rect 129 -155 161 -154
<< metal4 >>
rect 120 257 170 261
rect 120 225 129 257
rect 161 225 170 257
rect 120 221 170 225
rect 130 166 160 221
rect 120 162 170 166
rect 120 130 129 162
rect 161 130 170 162
rect 120 126 170 130
rect 130 71 160 126
rect 120 67 170 71
rect 120 35 129 67
rect 161 35 170 67
rect 120 31 170 35
rect 130 -24 160 31
rect 120 -28 170 -24
rect 120 -60 129 -28
rect 161 -60 170 -28
rect 120 -64 170 -60
rect 130 -119 160 -64
rect 120 -123 170 -119
rect 120 -155 129 -123
rect 161 -155 170 -123
rect 120 -159 170 -155
rect 130 -214 160 -159
rect 120 -254 170 -214
rect 130 -309 160 -254
rect 120 -349 170 -309
rect 130 -404 160 -349
rect 120 -444 170 -404
rect 130 -499 160 -444
rect 120 -539 170 -499
rect 130 -594 160 -539
rect 120 -634 170 -594
rect 130 -1934 160 -634
<< labels >>
rlabel metal1 -30 -724 -30 -724 7 VP
rlabel metal1 -30 -1379 -30 -1379 7 VN
rlabel metal1 54 351 54 351 1 col
rlabel metal1 -30 -234 -30 -234 3 Vgpc
rlabel metal1 -30 -664 -30 -664 3 Vc+
rlabel metal1 -30 -1224 -30 -1224 3 Vc-
rlabel metal1 -30 -1179 -30 -1179 3 Vgnc
rlabel metal1 -30 -1530 -30 -1530 3 Vref
rlabel metal3 145 -1930 145 -1930 1 SWref
rlabel metal2 150 -1930 150 -1930 1 SWc-
rlabel metal4 138 -1930 138 -1930 1 SWc+
<< end >>
